magic
tech sky130A
magscale 1 2
timestamp 1756452546
<< checkpaint >>
rect -3932 -3932 31903 34047
<< viali >>
rect 9781 27557 9815 27591
rect 10425 27557 10459 27591
rect 11069 27557 11103 27591
rect 11713 27557 11747 27591
rect 12357 27557 12391 27591
rect 14289 27557 14323 27591
rect 17509 27557 17543 27591
rect 20085 27557 20119 27591
rect 20729 27489 20763 27523
rect 9965 27421 9999 27455
rect 10609 27421 10643 27455
rect 11253 27421 11287 27455
rect 11897 27421 11931 27455
rect 12541 27421 12575 27455
rect 14473 27421 14507 27455
rect 17693 27421 17727 27455
rect 19441 27421 19475 27455
rect 19625 27421 19659 27455
rect 19717 27421 19751 27455
rect 20269 27421 20303 27455
rect 21373 27421 21407 27455
rect 21465 27421 21499 27455
rect 19257 27285 19291 27319
rect 21649 27285 21683 27319
rect 7941 27081 7975 27115
rect 10977 27013 11011 27047
rect 13737 27013 13771 27047
rect 14473 27013 14507 27047
rect 4997 26945 5031 26979
rect 7849 26945 7883 26979
rect 8309 26945 8343 26979
rect 9781 26945 9815 26979
rect 9965 26945 9999 26979
rect 10057 26945 10091 26979
rect 10241 26945 10275 26979
rect 10333 26945 10367 26979
rect 10425 26945 10459 26979
rect 10701 26945 10735 26979
rect 10885 26945 10919 26979
rect 11069 26945 11103 26979
rect 13001 26945 13035 26979
rect 13553 26945 13587 26979
rect 13645 26945 13679 26979
rect 13921 26945 13955 26979
rect 14289 26945 14323 26979
rect 14749 26945 14783 26979
rect 15117 26945 15151 26979
rect 16313 26945 16347 26979
rect 17109 26945 17143 26979
rect 17233 26945 17267 26979
rect 17325 26945 17359 26979
rect 17785 26945 17819 26979
rect 19053 26945 19087 26979
rect 20269 26945 20303 26979
rect 8401 26877 8435 26911
rect 8585 26877 8619 26911
rect 9505 26877 9539 26911
rect 14013 26877 14047 26911
rect 17877 26877 17911 26911
rect 17969 26877 18003 26911
rect 18797 26877 18831 26911
rect 16865 26809 16899 26843
rect 4813 26741 4847 26775
rect 7665 26741 7699 26775
rect 9597 26741 9631 26775
rect 10609 26741 10643 26775
rect 11253 26741 11287 26775
rect 12817 26741 12851 26775
rect 13369 26741 13403 26775
rect 14105 26741 14139 26775
rect 14657 26741 14691 26775
rect 14933 26741 14967 26775
rect 16405 26741 16439 26775
rect 17417 26741 17451 26775
rect 20177 26741 20211 26775
rect 20361 26741 20395 26775
rect 5825 26537 5859 26571
rect 8769 26537 8803 26571
rect 11897 26537 11931 26571
rect 8953 26469 8987 26503
rect 17601 26469 17635 26503
rect 7389 26401 7423 26435
rect 9505 26401 9539 26435
rect 10149 26401 10183 26435
rect 17509 26401 17543 26435
rect 19257 26401 19291 26435
rect 21005 26401 21039 26435
rect 4077 26333 4111 26367
rect 4445 26333 4479 26367
rect 7297 26333 7331 26367
rect 7656 26333 7690 26367
rect 12173 26333 12207 26367
rect 12449 26333 12483 26367
rect 12716 26333 12750 26367
rect 14289 26333 14323 26367
rect 15761 26333 15795 26367
rect 18981 26333 19015 26367
rect 21097 26333 21131 26367
rect 21281 26333 21315 26367
rect 23213 26333 23247 26367
rect 4712 26265 4746 26299
rect 10425 26265 10459 26299
rect 12081 26265 12115 26299
rect 14556 26265 14590 26299
rect 16037 26265 16071 26299
rect 18714 26265 18748 26299
rect 19533 26265 19567 26299
rect 23305 26265 23339 26299
rect 3893 26197 3927 26231
rect 7113 26197 7147 26231
rect 9321 26197 9355 26231
rect 9413 26197 9447 26231
rect 13829 26197 13863 26231
rect 15669 26197 15703 26231
rect 21189 26197 21223 26231
rect 5089 25993 5123 26027
rect 8401 25993 8435 26027
rect 9597 25993 9631 26027
rect 17141 25993 17175 26027
rect 18061 25993 18095 26027
rect 18797 25993 18831 26027
rect 18889 25993 18923 26027
rect 19257 25993 19291 26027
rect 5549 25925 5583 25959
rect 7266 25925 7300 25959
rect 11069 25925 11103 25959
rect 13277 25925 13311 25959
rect 15200 25925 15234 25959
rect 17785 25925 17819 25959
rect 21925 25925 21959 25959
rect 3617 25857 3651 25891
rect 3873 25857 3907 25891
rect 5457 25857 5491 25891
rect 6101 25857 6135 25891
rect 7021 25857 7055 25891
rect 9045 25857 9079 25891
rect 9321 25857 9355 25891
rect 11713 25857 11747 25891
rect 17049 25857 17083 25891
rect 17509 25857 17543 25891
rect 17693 25857 17727 25891
rect 17877 25857 17911 25891
rect 18613 25857 18647 25891
rect 22017 25857 22051 25891
rect 5641 25789 5675 25823
rect 11345 25789 11379 25823
rect 13001 25789 13035 25823
rect 14933 25789 14967 25823
rect 17233 25789 17267 25823
rect 19349 25789 19383 25823
rect 19441 25789 19475 25823
rect 21373 25789 21407 25823
rect 21649 25789 21683 25823
rect 22201 25789 22235 25823
rect 22477 25789 22511 25823
rect 24225 25789 24259 25823
rect 11621 25721 11655 25755
rect 14749 25721 14783 25755
rect 16681 25721 16715 25755
rect 4997 25653 5031 25687
rect 5917 25653 5951 25687
rect 9137 25653 9171 25687
rect 9505 25653 9539 25687
rect 16313 25653 16347 25687
rect 19901 25653 19935 25687
rect 4077 25449 4111 25483
rect 13001 25449 13035 25483
rect 15301 25449 15335 25483
rect 17417 25449 17451 25483
rect 19809 25449 19843 25483
rect 8769 25381 8803 25415
rect 22109 25381 22143 25415
rect 4721 25313 4755 25347
rect 7389 25313 7423 25347
rect 9597 25313 9631 25347
rect 13645 25313 13679 25347
rect 16129 25313 16163 25347
rect 21649 25313 21683 25347
rect 5365 25245 5399 25279
rect 5632 25245 5666 25279
rect 9137 25245 9171 25279
rect 9689 25245 9723 25279
rect 9873 25245 9907 25279
rect 10241 25245 10275 25279
rect 12265 25245 12299 25279
rect 13369 25245 13403 25279
rect 15485 25245 15519 25279
rect 17233 25245 17267 25279
rect 19257 25245 19291 25279
rect 19625 25245 19659 25279
rect 21097 25245 21131 25279
rect 21741 25245 21775 25279
rect 22937 25245 22971 25279
rect 4445 25177 4479 25211
rect 7656 25177 7690 25211
rect 10517 25177 10551 25211
rect 12173 25177 12207 25211
rect 15945 25177 15979 25211
rect 19441 25177 19475 25211
rect 19533 25177 19567 25211
rect 20821 25177 20855 25211
rect 4537 25109 4571 25143
rect 6745 25109 6779 25143
rect 8953 25109 8987 25143
rect 10057 25109 10091 25143
rect 11989 25109 12023 25143
rect 13461 25109 13495 25143
rect 15577 25109 15611 25143
rect 16037 25109 16071 25143
rect 23029 25109 23063 25143
rect 6377 24905 6411 24939
rect 8861 24905 8895 24939
rect 9229 24905 9263 24939
rect 10885 24905 10919 24939
rect 6745 24837 6779 24871
rect 6837 24837 6871 24871
rect 2513 24769 2547 24803
rect 3065 24769 3099 24803
rect 5457 24769 5491 24803
rect 8769 24769 8803 24803
rect 10333 24769 10367 24803
rect 10517 24769 10551 24803
rect 10609 24769 10643 24803
rect 10701 24769 10735 24803
rect 19165 24769 19199 24803
rect 19809 24769 19843 24803
rect 3157 24701 3191 24735
rect 3341 24701 3375 24735
rect 7021 24701 7055 24735
rect 8677 24701 8711 24735
rect 19901 24701 19935 24735
rect 20177 24701 20211 24735
rect 2697 24633 2731 24667
rect 2329 24565 2363 24599
rect 5273 24565 5307 24599
rect 19441 24565 19475 24599
rect 23857 24225 23891 24259
rect 1869 24157 1903 24191
rect 2136 24157 2170 24191
rect 4813 24157 4847 24191
rect 4905 24157 4939 24191
rect 13369 24157 13403 24191
rect 19901 24157 19935 24191
rect 20085 24157 20119 24191
rect 20177 24157 20211 24191
rect 22201 24157 22235 24191
rect 24409 24157 24443 24191
rect 5172 24089 5206 24123
rect 19993 24089 20027 24123
rect 20453 24089 20487 24123
rect 22109 24089 22143 24123
rect 23765 24089 23799 24123
rect 3249 24021 3283 24055
rect 4629 24021 4663 24055
rect 6285 24021 6319 24055
rect 13185 24021 13219 24055
rect 21925 24021 21959 24055
rect 23305 24021 23339 24055
rect 23673 24021 23707 24055
rect 24501 24021 24535 24055
rect 3525 23817 3559 23851
rect 3985 23817 4019 23851
rect 6377 23817 6411 23851
rect 6837 23817 6871 23851
rect 14841 23817 14875 23851
rect 20269 23817 20303 23851
rect 23397 23817 23431 23851
rect 4620 23749 4654 23783
rect 13154 23749 13188 23783
rect 19165 23749 19199 23783
rect 19349 23749 19383 23783
rect 23765 23749 23799 23783
rect 1777 23681 1811 23715
rect 2053 23681 2087 23715
rect 2309 23681 2343 23715
rect 3893 23681 3927 23715
rect 4353 23681 4387 23715
rect 6745 23681 6779 23715
rect 7941 23681 7975 23715
rect 11345 23681 11379 23715
rect 12633 23681 12667 23715
rect 14749 23681 14783 23715
rect 16129 23681 16163 23715
rect 16681 23681 16715 23715
rect 19533 23681 19567 23715
rect 19625 23681 19659 23715
rect 19809 23681 19843 23715
rect 19901 23681 19935 23715
rect 20177 23681 20211 23715
rect 20361 23681 20395 23715
rect 22477 23681 22511 23715
rect 23213 23681 23247 23715
rect 4169 23613 4203 23647
rect 7021 23613 7055 23647
rect 7665 23613 7699 23647
rect 7849 23613 7883 23647
rect 12909 23613 12943 23647
rect 15025 23613 15059 23647
rect 16037 23613 16071 23647
rect 16957 23613 16991 23647
rect 18705 23613 18739 23647
rect 20085 23613 20119 23647
rect 22385 23613 22419 23647
rect 22845 23613 22879 23647
rect 23489 23613 23523 23647
rect 1961 23545 1995 23579
rect 3433 23545 3467 23579
rect 5733 23545 5767 23579
rect 12817 23545 12851 23579
rect 14381 23545 14415 23579
rect 16497 23545 16531 23579
rect 8309 23477 8343 23511
rect 11253 23477 11287 23511
rect 14289 23477 14323 23511
rect 18889 23477 18923 23511
rect 19349 23477 19383 23511
rect 25237 23477 25271 23511
rect 5457 23273 5491 23307
rect 7113 23273 7147 23307
rect 12173 23273 12207 23307
rect 20177 23273 20211 23307
rect 20361 23273 20395 23307
rect 20085 23205 20119 23239
rect 1961 23137 1995 23171
rect 5917 23137 5951 23171
rect 6009 23137 6043 23171
rect 10425 23137 10459 23171
rect 12541 23137 12575 23171
rect 16681 23137 16715 23171
rect 18705 23137 18739 23171
rect 19625 23137 19659 23171
rect 19717 23137 19751 23171
rect 22477 23137 22511 23171
rect 4813 23069 4847 23103
rect 5089 23069 5123 23103
rect 5181 23069 5215 23103
rect 5825 23069 5859 23103
rect 6285 23069 6319 23103
rect 6561 23069 6595 23103
rect 6653 23069 6687 23103
rect 8493 23069 8527 23103
rect 8769 23069 8803 23103
rect 9781 23069 9815 23103
rect 10149 23069 10183 23103
rect 12449 23069 12483 23103
rect 12808 23069 12842 23103
rect 14105 23069 14139 23103
rect 15945 23069 15979 23103
rect 16093 23069 16127 23103
rect 16313 23069 16347 23103
rect 16451 23069 16485 23103
rect 18521 23069 18555 23103
rect 19257 23069 19291 23103
rect 19441 23069 19475 23103
rect 19809 23069 19843 23103
rect 19901 23069 19935 23103
rect 20729 23069 20763 23103
rect 20821 23069 20855 23103
rect 21189 23069 21223 23103
rect 22201 23069 22235 23103
rect 24409 23069 24443 23103
rect 24685 23069 24719 23103
rect 2228 23001 2262 23035
rect 4997 23001 5031 23035
rect 6469 23001 6503 23035
rect 8248 23001 8282 23035
rect 9965 23001 9999 23035
rect 10057 23001 10091 23035
rect 10701 23001 10735 23035
rect 12357 23001 12391 23035
rect 14372 23001 14406 23035
rect 16221 23001 16255 23035
rect 18429 23001 18463 23035
rect 20545 23001 20579 23035
rect 22753 23001 22787 23035
rect 24777 23001 24811 23035
rect 3341 22933 3375 22967
rect 5365 22933 5399 22967
rect 6837 22933 6871 22967
rect 8585 22933 8619 22967
rect 10333 22933 10367 22967
rect 13921 22933 13955 22967
rect 15485 22933 15519 22967
rect 16589 22933 16623 22967
rect 19349 22933 19383 22967
rect 20345 22933 20379 22967
rect 21005 22933 21039 22967
rect 22385 22933 22419 22967
rect 24225 22933 24259 22967
rect 24501 22933 24535 22967
rect 2329 22729 2363 22763
rect 2789 22729 2823 22763
rect 3157 22729 3191 22763
rect 6561 22729 6595 22763
rect 9505 22729 9539 22763
rect 11529 22729 11563 22763
rect 13369 22729 13403 22763
rect 13737 22729 13771 22763
rect 14381 22729 14415 22763
rect 14657 22729 14691 22763
rect 15025 22729 15059 22763
rect 22753 22729 22787 22763
rect 3249 22661 3283 22695
rect 3801 22661 3835 22695
rect 6898 22661 6932 22695
rect 8309 22661 8343 22695
rect 11805 22661 11839 22695
rect 12909 22661 12943 22695
rect 13001 22661 13035 22695
rect 15117 22661 15151 22695
rect 16681 22661 16715 22695
rect 17509 22661 17543 22695
rect 19441 22661 19475 22695
rect 22385 22661 22419 22695
rect 2513 22593 2547 22627
rect 3617 22593 3651 22627
rect 3893 22593 3927 22627
rect 3985 22593 4019 22627
rect 6377 22593 6411 22627
rect 8125 22593 8159 22627
rect 8401 22593 8435 22627
rect 8493 22593 8527 22627
rect 9321 22593 9355 22627
rect 9597 22593 9631 22627
rect 11713 22593 11747 22627
rect 11897 22593 11931 22627
rect 12081 22593 12115 22627
rect 12173 22593 12207 22627
rect 12357 22593 12391 22627
rect 12725 22593 12759 22627
rect 13093 22593 13127 22627
rect 13829 22593 13863 22627
rect 14565 22593 14599 22627
rect 17417 22593 17451 22627
rect 19717 22593 19751 22627
rect 20269 22593 20303 22627
rect 20545 22593 20579 22627
rect 20821 22593 20855 22627
rect 21373 22593 21407 22627
rect 23673 22593 23707 22627
rect 26341 22593 26375 22627
rect 3433 22525 3467 22559
rect 6653 22525 6687 22559
rect 9045 22525 9079 22559
rect 9873 22525 9907 22559
rect 11345 22525 11379 22559
rect 12633 22525 12667 22559
rect 14013 22525 14047 22559
rect 15209 22525 15243 22559
rect 17693 22525 17727 22559
rect 20085 22525 20119 22559
rect 22201 22525 22235 22559
rect 22293 22525 22327 22559
rect 23949 22525 23983 22559
rect 20453 22457 20487 22491
rect 21281 22457 21315 22491
rect 26525 22457 26559 22491
rect 4169 22389 4203 22423
rect 8033 22389 8067 22423
rect 8677 22389 8711 22423
rect 9137 22389 9171 22423
rect 12541 22389 12575 22423
rect 13277 22389 13311 22423
rect 25421 22389 25455 22423
rect 7205 22185 7239 22219
rect 12449 22185 12483 22219
rect 15761 22185 15795 22219
rect 21373 22185 21407 22219
rect 24041 22185 24075 22219
rect 21925 22117 21959 22151
rect 7849 22049 7883 22083
rect 8953 22049 8987 22083
rect 18153 22049 18187 22083
rect 21189 22049 21223 22083
rect 22109 22049 22143 22083
rect 23397 22049 23431 22083
rect 24501 22049 24535 22083
rect 2697 21981 2731 22015
rect 4905 21981 4939 22015
rect 5181 21981 5215 22015
rect 5365 21981 5399 22015
rect 7573 21981 7607 22015
rect 8585 21981 8619 22015
rect 11069 21981 11103 22015
rect 15209 21981 15243 22015
rect 15577 21981 15611 22015
rect 16313 21981 16347 22015
rect 16865 21981 16899 22015
rect 17417 21981 17451 22015
rect 17785 21981 17819 22015
rect 18521 21981 18555 22015
rect 19073 21981 19107 22015
rect 19809 21981 19843 22015
rect 19901 21981 19935 22015
rect 20361 21981 20395 22015
rect 20545 21981 20579 22015
rect 20637 21981 20671 22015
rect 21097 21981 21131 22015
rect 21557 21981 21591 22015
rect 21741 21981 21775 22015
rect 22017 21981 22051 22015
rect 22201 21981 22235 22015
rect 24225 21981 24259 22015
rect 24409 21981 24443 22015
rect 9198 21913 9232 21947
rect 11314 21913 11348 21947
rect 15393 21913 15427 21947
rect 15485 21913 15519 21947
rect 18061 21913 18095 21947
rect 18613 21913 18647 21947
rect 19349 21913 19383 21947
rect 19441 21913 19475 21947
rect 23581 21913 23615 21947
rect 2513 21845 2547 21879
rect 4721 21845 4755 21879
rect 5549 21845 5583 21879
rect 7665 21845 7699 21879
rect 8769 21845 8803 21879
rect 10333 21845 10367 21879
rect 16497 21845 16531 21879
rect 20821 21845 20855 21879
rect 23489 21845 23523 21879
rect 23949 21845 23983 21879
rect 7021 21641 7055 21675
rect 9137 21641 9171 21675
rect 9505 21641 9539 21675
rect 11161 21641 11195 21675
rect 11529 21641 11563 21675
rect 11897 21641 11931 21675
rect 15577 21641 15611 21675
rect 16037 21641 16071 21675
rect 21281 21641 21315 21675
rect 4528 21573 4562 21607
rect 6193 21573 6227 21607
rect 6745 21573 6779 21607
rect 19809 21573 19843 21607
rect 2053 21505 2087 21539
rect 2320 21505 2354 21539
rect 4261 21505 4295 21539
rect 5917 21505 5951 21539
rect 6377 21505 6411 21539
rect 6470 21505 6504 21539
rect 6653 21505 6687 21539
rect 6842 21505 6876 21539
rect 11345 21505 11379 21539
rect 11989 21505 12023 21539
rect 14197 21505 14231 21539
rect 14464 21505 14498 21539
rect 16129 21505 16163 21539
rect 19993 21505 20027 21539
rect 20361 21505 20395 21539
rect 20637 21505 20671 21539
rect 21189 21505 21223 21539
rect 22017 21505 22051 21539
rect 24317 21505 24351 21539
rect 25145 21505 25179 21539
rect 25789 21505 25823 21539
rect 6009 21437 6043 21471
rect 9597 21437 9631 21471
rect 9689 21437 9723 21471
rect 12081 21437 12115 21471
rect 16221 21437 16255 21471
rect 20545 21437 20579 21471
rect 21005 21437 21039 21471
rect 18521 21369 18555 21403
rect 3433 21301 3467 21335
rect 5641 21301 5675 21335
rect 5733 21301 5767 21335
rect 6193 21301 6227 21335
rect 15669 21301 15703 21335
rect 21925 21301 21959 21335
rect 24409 21301 24443 21335
rect 24777 21301 24811 21335
rect 25053 21301 25087 21335
rect 25697 21301 25731 21335
rect 3801 21097 3835 21131
rect 10057 21097 10091 21131
rect 14565 21097 14599 21131
rect 24777 21097 24811 21131
rect 1961 20961 1995 20995
rect 4445 20961 4479 20995
rect 5273 20961 5307 20995
rect 6469 20961 6503 20995
rect 22017 20961 22051 20995
rect 26525 20961 26559 20995
rect 4169 20893 4203 20927
rect 9505 20893 9539 20927
rect 9597 20893 9631 20927
rect 9781 20893 9815 20927
rect 9873 20893 9907 20927
rect 14749 20893 14783 20927
rect 16957 20893 16991 20927
rect 17141 20893 17175 20927
rect 17601 20893 17635 20927
rect 18337 20893 18371 20927
rect 18613 20893 18647 20927
rect 19349 20893 19383 20927
rect 19809 20893 19843 20927
rect 19901 20893 19935 20927
rect 20269 20893 20303 20927
rect 22109 20893 22143 20927
rect 23581 20893 23615 20927
rect 23949 20893 23983 20927
rect 24593 20893 24627 20927
rect 24685 20893 24719 20927
rect 2228 20825 2262 20859
rect 6009 20825 6043 20859
rect 6736 20825 6770 20859
rect 19441 20825 19475 20859
rect 19993 20825 20027 20859
rect 23765 20825 23799 20859
rect 23857 20825 23891 20859
rect 26249 20825 26283 20859
rect 3341 20757 3375 20791
rect 4261 20757 4295 20791
rect 7849 20757 7883 20791
rect 16773 20757 16807 20791
rect 18889 20757 18923 20791
rect 22201 20757 22235 20791
rect 24133 20757 24167 20791
rect 2421 20553 2455 20587
rect 2881 20553 2915 20587
rect 3249 20553 3283 20587
rect 4905 20553 4939 20587
rect 5273 20553 5307 20587
rect 6745 20553 6779 20587
rect 7021 20553 7055 20587
rect 7389 20553 7423 20587
rect 21097 20553 21131 20587
rect 21465 20553 21499 20587
rect 24041 20553 24075 20587
rect 24777 20553 24811 20587
rect 25145 20553 25179 20587
rect 4077 20485 4111 20519
rect 5365 20485 5399 20519
rect 7481 20485 7515 20519
rect 9965 20485 9999 20519
rect 14105 20485 14139 20519
rect 17417 20485 17451 20519
rect 17969 20485 18003 20519
rect 18797 20485 18831 20519
rect 20453 20485 20487 20519
rect 24133 20485 24167 20519
rect 2605 20417 2639 20451
rect 3801 20417 3835 20451
rect 3985 20417 4019 20451
rect 4169 20417 4203 20451
rect 6929 20417 6963 20451
rect 9873 20417 9907 20451
rect 13277 20417 13311 20451
rect 13553 20417 13587 20451
rect 13829 20417 13863 20451
rect 13977 20417 14011 20451
rect 14197 20417 14231 20451
rect 14335 20417 14369 20451
rect 17509 20417 17543 20451
rect 18705 20417 18739 20451
rect 19441 20417 19475 20451
rect 19901 20417 19935 20451
rect 19993 20417 20027 20451
rect 20269 20417 20303 20451
rect 21833 20417 21867 20451
rect 22661 20417 22695 20451
rect 23581 20417 23615 20451
rect 25053 20417 25087 20451
rect 25513 20417 25547 20451
rect 26065 20417 26099 20451
rect 3341 20349 3375 20383
rect 3525 20349 3559 20383
rect 5457 20349 5491 20383
rect 7573 20349 7607 20383
rect 10149 20349 10183 20383
rect 16957 20349 16991 20383
rect 17877 20349 17911 20383
rect 18245 20349 18279 20383
rect 18337 20349 18371 20383
rect 19257 20349 19291 20383
rect 19533 20349 19567 20383
rect 20913 20349 20947 20383
rect 21005 20349 21039 20383
rect 22477 20349 22511 20383
rect 24501 20349 24535 20383
rect 25237 20349 25271 20383
rect 25421 20349 25455 20383
rect 4353 20281 4387 20315
rect 24298 20281 24332 20315
rect 24961 20281 24995 20315
rect 25605 20281 25639 20315
rect 9505 20213 9539 20247
rect 13093 20213 13127 20247
rect 13369 20213 13403 20247
rect 14473 20213 14507 20247
rect 20545 20213 20579 20247
rect 22017 20213 22051 20247
rect 23673 20213 23707 20247
rect 24409 20213 24443 20247
rect 25789 20213 25823 20247
rect 14105 20009 14139 20043
rect 19257 20009 19291 20043
rect 24041 20009 24075 20043
rect 24685 20009 24719 20043
rect 3341 19941 3375 19975
rect 22937 19941 22971 19975
rect 8953 19873 8987 19907
rect 14657 19873 14691 19907
rect 18061 19873 18095 19907
rect 22017 19873 22051 19907
rect 22477 19873 22511 19907
rect 1961 19805 1995 19839
rect 3801 19805 3835 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 4169 19805 4203 19839
rect 4721 19805 4755 19839
rect 6745 19805 6779 19839
rect 8585 19805 8619 19839
rect 10609 19805 10643 19839
rect 11069 19805 11103 19839
rect 12541 19805 12575 19839
rect 12808 19805 12842 19839
rect 14473 19805 14507 19839
rect 16313 19805 16347 19839
rect 17049 19805 17083 19839
rect 17417 19805 17451 19839
rect 17785 19805 17819 19839
rect 18521 19805 18555 19839
rect 19073 19805 19107 19839
rect 19533 19805 19567 19839
rect 19809 19805 19843 19839
rect 20085 19805 20119 19839
rect 22293 19805 22327 19839
rect 22569 19805 22603 19839
rect 23949 19805 23983 19839
rect 24869 19805 24903 19839
rect 24961 19805 24995 19839
rect 25237 19805 25271 19839
rect 25513 19805 25547 19839
rect 2228 19737 2262 19771
rect 6990 19737 7024 19771
rect 9198 19737 9232 19771
rect 11336 19737 11370 19771
rect 14565 19737 14599 19771
rect 18153 19737 18187 19771
rect 18613 19737 18647 19771
rect 25053 19737 25087 19771
rect 25421 19737 25455 19771
rect 4353 19669 4387 19703
rect 8125 19669 8159 19703
rect 8769 19669 8803 19703
rect 10333 19669 10367 19703
rect 12449 19669 12483 19703
rect 13921 19669 13955 19703
rect 16681 19669 16715 19703
rect 20545 19669 20579 19703
rect 2421 19465 2455 19499
rect 2789 19465 2823 19499
rect 3157 19465 3191 19499
rect 6561 19465 6595 19499
rect 7849 19465 7883 19499
rect 9413 19465 9447 19499
rect 11529 19465 11563 19499
rect 12265 19465 12299 19499
rect 14197 19465 14231 19499
rect 14565 19465 14599 19499
rect 14657 19465 14691 19499
rect 18613 19465 18647 19499
rect 20469 19465 20503 19499
rect 20637 19465 20671 19499
rect 21833 19465 21867 19499
rect 4721 19397 4755 19431
rect 7021 19397 7055 19431
rect 7113 19397 7147 19431
rect 10057 19397 10091 19431
rect 11161 19397 11195 19431
rect 12992 19397 13026 19431
rect 16773 19397 16807 19431
rect 20269 19397 20303 19431
rect 2605 19329 2639 19363
rect 3249 19329 3283 19363
rect 5457 19329 5491 19363
rect 6377 19329 6411 19363
rect 6745 19329 6779 19363
rect 6893 19329 6927 19363
rect 7210 19329 7244 19363
rect 7941 19329 7975 19363
rect 9505 19329 9539 19363
rect 9965 19329 9999 19363
rect 10425 19329 10459 19363
rect 11713 19329 11747 19363
rect 12173 19329 12207 19363
rect 12725 19329 12759 19363
rect 15945 19329 15979 19363
rect 16865 19329 16899 19363
rect 17233 19329 17267 19363
rect 17325 19329 17359 19363
rect 17785 19329 17819 19363
rect 18337 19329 18371 19363
rect 18981 19329 19015 19363
rect 19533 19329 19567 19363
rect 19717 19329 19751 19363
rect 3433 19261 3467 19295
rect 8125 19261 8159 19295
rect 9045 19261 9079 19295
rect 10241 19261 10275 19295
rect 12357 19261 12391 19295
rect 14749 19261 14783 19295
rect 23305 19261 23339 19295
rect 23581 19261 23615 19295
rect 7389 19193 7423 19227
rect 7481 19193 7515 19227
rect 9229 19193 9263 19227
rect 11805 19193 11839 19227
rect 14105 19193 14139 19227
rect 8769 19125 8803 19159
rect 9137 19125 9171 19159
rect 9597 19125 9631 19159
rect 20453 19125 20487 19159
rect 8493 18921 8527 18955
rect 11069 18921 11103 18955
rect 12173 18921 12207 18955
rect 22201 18921 22235 18955
rect 26433 18921 26467 18955
rect 4629 18785 4663 18819
rect 7573 18785 7607 18819
rect 14749 18785 14783 18819
rect 17601 18785 17635 18819
rect 19441 18785 19475 18819
rect 2329 18717 2363 18751
rect 3617 18717 3651 18751
rect 4813 18717 4847 18751
rect 4906 18717 4940 18751
rect 5278 18717 5312 18751
rect 6929 18717 6963 18751
rect 7389 18717 7423 18751
rect 7849 18717 7883 18751
rect 7942 18717 7976 18751
rect 8125 18717 8159 18751
rect 8355 18717 8389 18751
rect 9045 18717 9079 18751
rect 9505 18717 9539 18751
rect 9689 18717 9723 18751
rect 11621 18717 11655 18751
rect 11713 18717 11747 18751
rect 11897 18717 11931 18751
rect 11989 18717 12023 18751
rect 16589 18717 16623 18751
rect 18061 18717 18095 18751
rect 19257 18717 19291 18751
rect 22109 18717 22143 18751
rect 24685 18717 24719 18751
rect 4353 18649 4387 18683
rect 5089 18649 5123 18683
rect 5181 18649 5215 18683
rect 8217 18649 8251 18683
rect 9934 18649 9968 18683
rect 15016 18649 15050 18683
rect 17417 18649 17451 18683
rect 17693 18649 17727 18683
rect 18153 18649 18187 18683
rect 18245 18649 18279 18683
rect 24961 18649 24995 18683
rect 2145 18581 2179 18615
rect 3433 18581 3467 18615
rect 3985 18581 4019 18615
rect 4445 18581 4479 18615
rect 5457 18581 5491 18615
rect 6745 18581 6779 18615
rect 7021 18581 7055 18615
rect 7481 18581 7515 18615
rect 9229 18581 9263 18615
rect 9321 18581 9355 18615
rect 16129 18581 16163 18615
rect 3893 18377 3927 18411
rect 5365 18377 5399 18411
rect 5457 18377 5491 18411
rect 7849 18377 7883 18411
rect 8401 18377 8435 18411
rect 10333 18377 10367 18411
rect 15117 18377 15151 18411
rect 15761 18377 15795 18411
rect 25789 18377 25823 18411
rect 26249 18377 26283 18411
rect 4252 18309 4286 18343
rect 9220 18309 9254 18343
rect 11161 18309 11195 18343
rect 18337 18309 18371 18343
rect 18889 18309 18923 18343
rect 2053 18241 2087 18275
rect 2237 18241 2271 18275
rect 2513 18241 2547 18275
rect 2780 18241 2814 18275
rect 3985 18241 4019 18275
rect 5641 18241 5675 18275
rect 6009 18241 6043 18275
rect 6469 18241 6503 18275
rect 6725 18241 6759 18275
rect 8309 18241 8343 18275
rect 8953 18241 8987 18275
rect 10425 18241 10459 18275
rect 15301 18241 15335 18275
rect 16129 18241 16163 18275
rect 17601 18241 17635 18275
rect 18245 18241 18279 18275
rect 18429 18241 18463 18275
rect 22201 18241 22235 18275
rect 24041 18241 24075 18275
rect 26065 18241 26099 18275
rect 26157 18241 26191 18275
rect 1409 18173 1443 18207
rect 8585 18173 8619 18207
rect 16221 18173 16255 18207
rect 16405 18173 16439 18207
rect 16773 18173 16807 18207
rect 18797 18173 18831 18207
rect 22477 18173 22511 18207
rect 24317 18173 24351 18207
rect 6193 18105 6227 18139
rect 2329 18037 2363 18071
rect 7941 18037 7975 18071
rect 23949 18037 23983 18071
rect 25973 18037 26007 18071
rect 3801 17833 3835 17867
rect 5365 17833 5399 17867
rect 8033 17833 8067 17867
rect 9413 17833 9447 17867
rect 10425 17833 10459 17867
rect 23397 17833 23431 17867
rect 23857 17833 23891 17867
rect 24133 17833 24167 17867
rect 26157 17833 26191 17867
rect 2881 17765 2915 17799
rect 4353 17697 4387 17731
rect 4813 17697 4847 17731
rect 6653 17697 6687 17731
rect 10057 17697 10091 17731
rect 12449 17697 12483 17731
rect 12633 17697 12667 17731
rect 18613 17697 18647 17731
rect 21649 17697 21683 17731
rect 21925 17697 21959 17731
rect 24409 17697 24443 17731
rect 1501 17629 1535 17663
rect 1768 17629 1802 17663
rect 4169 17629 4203 17663
rect 4997 17629 5031 17663
rect 6920 17629 6954 17663
rect 9781 17629 9815 17663
rect 10609 17629 10643 17663
rect 10977 17629 11011 17663
rect 12357 17629 12391 17663
rect 16037 17629 16071 17663
rect 19257 17629 19291 17663
rect 23673 17629 23707 17663
rect 23949 17629 23983 17663
rect 24041 17629 24075 17663
rect 26249 17629 26283 17663
rect 4261 17561 4295 17595
rect 10701 17561 10735 17595
rect 10793 17561 10827 17595
rect 18337 17561 18371 17595
rect 23581 17561 23615 17595
rect 24685 17561 24719 17595
rect 26341 17561 26375 17595
rect 4905 17493 4939 17527
rect 9873 17493 9907 17527
rect 11989 17493 12023 17527
rect 17969 17493 18003 17527
rect 18429 17493 18463 17527
rect 19441 17493 19475 17527
rect 3065 17289 3099 17323
rect 13001 17289 13035 17323
rect 17693 17289 17727 17323
rect 19165 17289 19199 17323
rect 21833 17289 21867 17323
rect 24593 17289 24627 17323
rect 3525 17221 3559 17255
rect 12541 17221 12575 17255
rect 18030 17221 18064 17255
rect 20370 17221 20404 17255
rect 23305 17221 23339 17255
rect 1685 17153 1719 17187
rect 1952 17153 1986 17187
rect 4169 17153 4203 17187
rect 9781 17153 9815 17187
rect 10517 17153 10551 17187
rect 13185 17153 13219 17187
rect 13277 17153 13311 17187
rect 13461 17153 13495 17187
rect 13553 17153 13587 17187
rect 14289 17153 14323 17187
rect 14556 17153 14590 17187
rect 15761 17153 15795 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 16129 17153 16163 17187
rect 17509 17153 17543 17187
rect 21649 17153 21683 17187
rect 3617 17085 3651 17119
rect 3709 17085 3743 17119
rect 12633 17085 12667 17119
rect 12817 17085 12851 17119
rect 17785 17085 17819 17119
rect 20637 17085 20671 17119
rect 23581 17085 23615 17119
rect 26065 17085 26099 17119
rect 26341 17085 26375 17119
rect 3157 17017 3191 17051
rect 4353 16949 4387 16983
rect 10333 16949 10367 16983
rect 12173 16949 12207 16983
rect 15669 16949 15703 16983
rect 16313 16949 16347 16983
rect 19257 16949 19291 16983
rect 21557 16949 21591 16983
rect 2237 16745 2271 16779
rect 4905 16745 4939 16779
rect 11069 16745 11103 16779
rect 13185 16745 13219 16779
rect 13829 16745 13863 16779
rect 19257 16745 19291 16779
rect 20085 16745 20119 16779
rect 6745 16609 6779 16643
rect 6837 16609 6871 16643
rect 9689 16609 9723 16643
rect 11805 16609 11839 16643
rect 15025 16609 15059 16643
rect 15301 16609 15335 16643
rect 17325 16609 17359 16643
rect 17693 16609 17727 16643
rect 19901 16609 19935 16643
rect 20177 16609 20211 16643
rect 20729 16609 20763 16643
rect 21005 16609 21039 16643
rect 2421 16541 2455 16575
rect 4261 16541 4295 16575
rect 4354 16541 4388 16575
rect 4629 16541 4663 16575
rect 4767 16541 4801 16575
rect 6653 16541 6687 16575
rect 7113 16541 7147 16575
rect 7481 16541 7515 16575
rect 9956 16541 9990 16575
rect 11253 16541 11287 16575
rect 11529 16541 11563 16575
rect 13277 16541 13311 16575
rect 13461 16541 13495 16575
rect 13645 16541 13679 16575
rect 14197 16541 14231 16575
rect 17233 16541 17267 16575
rect 19625 16541 19659 16575
rect 20361 16541 20395 16575
rect 4537 16473 4571 16507
rect 7297 16473 7331 16507
rect 7389 16473 7423 16507
rect 12050 16473 12084 16507
rect 13553 16473 13587 16507
rect 14841 16473 14875 16507
rect 15568 16473 15602 16507
rect 17141 16473 17175 16507
rect 17960 16473 17994 16507
rect 20085 16473 20119 16507
rect 22569 16473 22603 16507
rect 23397 16473 23431 16507
rect 6285 16405 6319 16439
rect 7665 16405 7699 16439
rect 11437 16405 11471 16439
rect 11713 16405 11747 16439
rect 14381 16405 14415 16439
rect 14473 16405 14507 16439
rect 14933 16405 14967 16439
rect 16681 16405 16715 16439
rect 16773 16405 16807 16439
rect 19073 16405 19107 16439
rect 19717 16405 19751 16439
rect 20545 16405 20579 16439
rect 22477 16405 22511 16439
rect 2881 16201 2915 16235
rect 3433 16201 3467 16235
rect 7757 16201 7791 16235
rect 7941 16201 7975 16235
rect 9321 16201 9355 16235
rect 10241 16201 10275 16235
rect 10609 16201 10643 16235
rect 13645 16201 13679 16235
rect 14381 16201 14415 16235
rect 15945 16201 15979 16235
rect 17325 16201 17359 16235
rect 17877 16201 17911 16235
rect 18153 16201 18187 16235
rect 18521 16201 18555 16235
rect 19993 16201 20027 16235
rect 22937 16201 22971 16235
rect 14718 16133 14752 16167
rect 17049 16133 17083 16167
rect 21833 16133 21867 16167
rect 1501 16065 1535 16099
rect 1768 16065 1802 16099
rect 3341 16065 3375 16099
rect 3985 16065 4019 16099
rect 5917 16065 5951 16099
rect 6377 16065 6411 16099
rect 6633 16065 6667 16099
rect 8125 16065 8159 16099
rect 8401 16065 8435 16099
rect 9229 16065 9263 16099
rect 9689 16065 9723 16099
rect 11161 16065 11195 16099
rect 11969 16065 12003 16099
rect 13553 16065 13587 16099
rect 14197 16065 14231 16099
rect 16129 16065 16163 16099
rect 16681 16065 16715 16099
rect 16829 16065 16863 16099
rect 16957 16065 16991 16099
rect 17187 16065 17221 16099
rect 18061 16065 18095 16099
rect 18981 16065 19015 16099
rect 19073 16065 19107 16099
rect 19257 16065 19291 16099
rect 19349 16065 19383 16099
rect 19625 16065 19659 16099
rect 19809 16065 19843 16099
rect 21557 16065 21591 16099
rect 23029 16065 23063 16099
rect 26249 16065 26283 16099
rect 26341 16065 26375 16099
rect 3617 15997 3651 16031
rect 9781 15997 9815 16031
rect 9965 15997 9999 16031
rect 10701 15997 10735 16031
rect 10885 15997 10919 16031
rect 11713 15997 11747 16031
rect 13737 15997 13771 16031
rect 14473 15997 14507 16031
rect 18613 15997 18647 16031
rect 18705 15997 18739 16031
rect 22569 15997 22603 16031
rect 2973 15929 3007 15963
rect 6101 15929 6135 15963
rect 11345 15929 11379 15963
rect 15853 15929 15887 15963
rect 19533 15929 19567 15963
rect 3801 15861 3835 15895
rect 8217 15861 8251 15895
rect 9045 15861 9079 15895
rect 13093 15861 13127 15895
rect 13185 15861 13219 15895
rect 26157 15861 26191 15895
rect 26433 15861 26467 15895
rect 3801 15657 3835 15691
rect 4629 15657 4663 15691
rect 6929 15657 6963 15691
rect 10333 15657 10367 15691
rect 13277 15657 13311 15691
rect 14841 15657 14875 15691
rect 18981 15657 19015 15691
rect 10425 15589 10459 15623
rect 19349 15589 19383 15623
rect 4445 15521 4479 15555
rect 5549 15521 5583 15555
rect 11897 15521 11931 15555
rect 15485 15521 15519 15555
rect 20729 15521 20763 15555
rect 2237 15453 2271 15487
rect 2504 15453 2538 15487
rect 4813 15453 4847 15487
rect 4997 15453 5031 15487
rect 5181 15453 5215 15487
rect 8134 15453 8168 15487
rect 8401 15453 8435 15487
rect 8953 15453 8987 15487
rect 10609 15453 10643 15487
rect 10701 15453 10735 15487
rect 10885 15453 10919 15487
rect 10977 15453 11011 15487
rect 12153 15453 12187 15487
rect 15209 15453 15243 15487
rect 18429 15453 18463 15487
rect 18705 15453 18739 15487
rect 18797 15453 18831 15487
rect 21833 15453 21867 15487
rect 23029 15453 23063 15487
rect 24409 15453 24443 15487
rect 26249 15453 26283 15487
rect 4905 15385 4939 15419
rect 5816 15385 5850 15419
rect 9198 15385 9232 15419
rect 18613 15385 18647 15419
rect 20462 15385 20496 15419
rect 24685 15385 24719 15419
rect 3617 15317 3651 15351
rect 4169 15317 4203 15351
rect 4261 15317 4295 15351
rect 7021 15317 7055 15351
rect 15301 15317 15335 15351
rect 22937 15317 22971 15351
rect 26157 15317 26191 15351
rect 26341 15317 26375 15351
rect 2145 15113 2179 15147
rect 4261 15113 4295 15147
rect 4721 15113 4755 15147
rect 5917 15113 5951 15147
rect 6745 15113 6779 15147
rect 7665 15113 7699 15147
rect 8125 15113 8159 15147
rect 9873 15113 9907 15147
rect 10517 15113 10551 15147
rect 19257 15113 19291 15147
rect 19349 15113 19383 15147
rect 19717 15113 19751 15147
rect 19993 15113 20027 15147
rect 3148 15045 3182 15079
rect 10149 15045 10183 15079
rect 10241 15045 10275 15079
rect 14013 15045 14047 15079
rect 2329 14977 2363 15011
rect 6101 14977 6135 15011
rect 7757 14977 7791 15011
rect 8217 14977 8251 15011
rect 8500 14977 8534 15011
rect 8760 14977 8794 15011
rect 9965 14977 9999 15011
rect 10333 14977 10367 15011
rect 19809 14977 19843 15011
rect 25053 14977 25087 15011
rect 2881 14909 2915 14943
rect 4813 14909 4847 14943
rect 4905 14909 4939 14943
rect 6837 14909 6871 14943
rect 6929 14909 6963 14943
rect 7481 14909 7515 14943
rect 19165 14909 19199 14943
rect 21833 14909 21867 14943
rect 22109 14909 22143 14943
rect 25605 14909 25639 14943
rect 25973 14909 26007 14943
rect 6377 14841 6411 14875
rect 8401 14841 8435 14875
rect 4353 14773 4387 14807
rect 15301 14773 15335 14807
rect 23581 14773 23615 14807
rect 25145 14773 25179 14807
rect 26525 14773 26559 14807
rect 3249 14569 3283 14603
rect 9045 14569 9079 14603
rect 16773 14569 16807 14603
rect 19349 14569 19383 14603
rect 26341 14569 26375 14603
rect 18337 14501 18371 14535
rect 9597 14433 9631 14467
rect 15117 14433 15151 14467
rect 21189 14433 21223 14467
rect 21465 14433 21499 14467
rect 24685 14433 24719 14467
rect 3433 14365 3467 14399
rect 9413 14365 9447 14399
rect 14473 14365 14507 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 15761 14365 15795 14399
rect 16221 14365 16255 14399
rect 16313 14365 16347 14399
rect 16497 14365 16531 14399
rect 16589 14365 16623 14399
rect 18475 14365 18509 14399
rect 18705 14365 18739 14399
rect 18888 14365 18922 14399
rect 18981 14365 19015 14399
rect 19533 14365 19567 14399
rect 23213 14365 23247 14399
rect 24409 14365 24443 14399
rect 26433 14365 26467 14399
rect 9505 14297 9539 14331
rect 14933 14297 14967 14331
rect 15577 14297 15611 14331
rect 18613 14297 18647 14331
rect 23121 14297 23155 14331
rect 14289 14229 14323 14263
rect 14565 14229 14599 14263
rect 15025 14229 15059 14263
rect 15945 14229 15979 14263
rect 22937 14229 22971 14263
rect 26157 14229 26191 14263
rect 13553 14025 13587 14059
rect 15025 14025 15059 14059
rect 16497 14025 16531 14059
rect 17049 14025 17083 14059
rect 18797 14025 18831 14059
rect 19257 14025 19291 14059
rect 13912 13957 13946 13991
rect 17877 13957 17911 13991
rect 22293 13957 22327 13991
rect 24225 13957 24259 13991
rect 10609 13889 10643 13923
rect 10701 13889 10735 13923
rect 10885 13889 10919 13923
rect 10987 13889 11021 13923
rect 11713 13889 11747 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 13369 13889 13403 13923
rect 15384 13889 15418 13923
rect 17141 13889 17175 13923
rect 17969 13889 18003 13923
rect 20370 13889 20404 13923
rect 24133 13889 24167 13923
rect 11529 13821 11563 13855
rect 13645 13821 13679 13855
rect 15117 13821 15151 13855
rect 17233 13821 17267 13855
rect 18061 13821 18095 13855
rect 18521 13821 18555 13855
rect 18705 13821 18739 13855
rect 20637 13821 20671 13855
rect 22017 13821 22051 13855
rect 23765 13821 23799 13855
rect 24409 13821 24443 13855
rect 10425 13753 10459 13787
rect 12357 13685 12391 13719
rect 16681 13685 16715 13719
rect 17509 13685 17543 13719
rect 19165 13685 19199 13719
rect 24672 13685 24706 13719
rect 26157 13685 26191 13719
rect 5917 13481 5951 13515
rect 11437 13481 11471 13515
rect 15485 13481 15519 13515
rect 15761 13481 15795 13515
rect 19073 13481 19107 13515
rect 23029 13481 23063 13515
rect 5273 13413 5307 13447
rect 6101 13413 6135 13447
rect 10885 13413 10919 13447
rect 19257 13413 19291 13447
rect 1961 13345 1995 13379
rect 4261 13345 4295 13379
rect 4445 13345 4479 13379
rect 5733 13345 5767 13379
rect 7205 13345 7239 13379
rect 9689 13345 9723 13379
rect 10241 13345 10275 13379
rect 12817 13345 12851 13379
rect 14105 13345 14139 13379
rect 17049 13345 17083 13379
rect 24777 13345 24811 13379
rect 25053 13345 25087 13379
rect 2237 13277 2271 13311
rect 2697 13277 2731 13311
rect 2973 13277 3007 13311
rect 4629 13277 4663 13311
rect 4722 13277 4756 13311
rect 4905 13277 4939 13311
rect 5094 13277 5128 13311
rect 5641 13277 5675 13311
rect 5917 13277 5951 13311
rect 6193 13277 6227 13311
rect 10517 13277 10551 13311
rect 10977 13277 11011 13311
rect 12550 13277 12584 13311
rect 13277 13277 13311 13311
rect 15945 13277 15979 13311
rect 16497 13277 16531 13311
rect 16957 13277 16991 13311
rect 18521 13277 18555 13311
rect 18889 13277 18923 13311
rect 20637 13277 20671 13311
rect 23121 13277 23155 13311
rect 4997 13209 5031 13243
rect 7021 13209 7055 13243
rect 9505 13209 9539 13243
rect 14350 13209 14384 13243
rect 17294 13209 17328 13243
rect 18705 13209 18739 13243
rect 18797 13209 18831 13243
rect 20370 13209 20404 13243
rect 2513 13141 2547 13175
rect 2789 13141 2823 13175
rect 3801 13141 3835 13175
rect 4169 13141 4203 13175
rect 6377 13141 6411 13175
rect 6561 13141 6595 13175
rect 6929 13141 6963 13175
rect 9137 13141 9171 13175
rect 9597 13141 9631 13175
rect 10425 13141 10459 13175
rect 11161 13141 11195 13175
rect 13093 13141 13127 13175
rect 16681 13141 16715 13175
rect 16773 13141 16807 13175
rect 18429 13141 18463 13175
rect 26525 13141 26559 13175
rect 2053 12937 2087 12971
rect 3801 12937 3835 12971
rect 4169 12937 4203 12971
rect 6193 12937 6227 12971
rect 7757 12937 7791 12971
rect 9965 12937 9999 12971
rect 11897 12937 11931 12971
rect 12265 12937 12299 12971
rect 14381 12937 14415 12971
rect 14749 12937 14783 12971
rect 18061 12937 18095 12971
rect 18153 12937 18187 12971
rect 18521 12937 18555 12971
rect 18613 12937 18647 12971
rect 19349 12937 19383 12971
rect 19441 12937 19475 12971
rect 19993 12937 20027 12971
rect 2596 12869 2630 12903
rect 4997 12869 5031 12903
rect 5825 12869 5859 12903
rect 6622 12869 6656 12903
rect 8125 12869 8159 12903
rect 12900 12869 12934 12903
rect 14841 12869 14875 12903
rect 16926 12869 16960 12903
rect 26065 12869 26099 12903
rect 1409 12801 1443 12835
rect 5089 12801 5123 12835
rect 8033 12801 8067 12835
rect 8217 12801 8251 12835
rect 8401 12801 8435 12835
rect 8749 12801 8783 12835
rect 11078 12801 11112 12835
rect 19809 12801 19843 12835
rect 22017 12801 22051 12835
rect 26341 12801 26375 12835
rect 2329 12733 2363 12767
rect 4261 12733 4295 12767
rect 4353 12733 4387 12767
rect 5273 12733 5307 12767
rect 5641 12733 5675 12767
rect 5733 12733 5767 12767
rect 6377 12733 6411 12767
rect 8493 12733 8527 12767
rect 11345 12733 11379 12767
rect 11621 12733 11655 12767
rect 11805 12733 11839 12767
rect 12633 12733 12667 12767
rect 14933 12733 14967 12767
rect 16681 12733 16715 12767
rect 18705 12733 18739 12767
rect 19533 12733 19567 12767
rect 3709 12665 3743 12699
rect 7849 12665 7883 12699
rect 4629 12597 4663 12631
rect 9873 12597 9907 12631
rect 14013 12597 14047 12631
rect 18981 12597 19015 12631
rect 21833 12597 21867 12631
rect 24593 12597 24627 12631
rect 3249 12393 3283 12427
rect 5549 12393 5583 12427
rect 7389 12393 7423 12427
rect 8585 12393 8619 12427
rect 13093 12393 13127 12427
rect 18981 12393 19015 12427
rect 22661 12393 22695 12427
rect 6009 12257 6043 12291
rect 9045 12257 9079 12291
rect 10977 12257 11011 12291
rect 11069 12257 11103 12291
rect 13737 12257 13771 12291
rect 20913 12257 20947 12291
rect 21189 12257 21223 12291
rect 24961 12257 24995 12291
rect 1869 12189 1903 12223
rect 4077 12189 4111 12223
rect 4169 12189 4203 12223
rect 8769 12189 8803 12223
rect 18797 12189 18831 12223
rect 20821 12189 20855 12223
rect 22937 12189 22971 12223
rect 23949 12189 23983 12223
rect 24777 12189 24811 12223
rect 25789 12189 25823 12223
rect 2136 12121 2170 12155
rect 4436 12121 4470 12155
rect 6276 12121 6310 12155
rect 9312 12121 9346 12155
rect 10885 12121 10919 12155
rect 13461 12121 13495 12155
rect 22845 12121 22879 12155
rect 3893 12053 3927 12087
rect 10425 12053 10459 12087
rect 10517 12053 10551 12087
rect 13553 12053 13587 12087
rect 20637 12053 20671 12087
rect 23765 12053 23799 12087
rect 24409 12053 24443 12087
rect 24869 12053 24903 12087
rect 25697 12053 25731 12087
rect 2973 11849 3007 11883
rect 4629 11849 4663 11883
rect 5917 11849 5951 11883
rect 6377 11849 6411 11883
rect 9413 11849 9447 11883
rect 10977 11849 11011 11883
rect 21649 11849 21683 11883
rect 22017 11849 22051 11883
rect 22385 11849 22419 11883
rect 10609 11781 10643 11815
rect 10701 11781 10735 11815
rect 20177 11781 20211 11815
rect 23673 11781 23707 11815
rect 25329 11781 25363 11815
rect 1593 11713 1627 11747
rect 1860 11713 1894 11747
rect 3433 11713 3467 11747
rect 4169 11713 4203 11747
rect 4353 11713 4387 11747
rect 4813 11713 4847 11747
rect 5641 11713 5675 11747
rect 5733 11713 5767 11747
rect 6561 11713 6595 11747
rect 9597 11713 9631 11747
rect 10425 11713 10459 11747
rect 10793 11713 10827 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 25421 11713 25455 11747
rect 25513 11713 25547 11747
rect 3525 11645 3559 11679
rect 3709 11645 3743 11679
rect 19901 11645 19935 11679
rect 22477 11645 22511 11679
rect 22569 11645 22603 11679
rect 23397 11645 23431 11679
rect 3065 11577 3099 11611
rect 25145 11577 25179 11611
rect 4537 11509 4571 11543
rect 14289 11509 14323 11543
rect 25605 11509 25639 11543
rect 2145 11305 2179 11339
rect 20821 11305 20855 11339
rect 21741 11305 21775 11339
rect 26157 11305 26191 11339
rect 12357 11237 12391 11271
rect 15485 11237 15519 11271
rect 18797 11237 18831 11271
rect 12909 11169 12943 11203
rect 15945 11169 15979 11203
rect 16129 11169 16163 11203
rect 18153 11169 18187 11203
rect 21373 11169 21407 11203
rect 24409 11169 24443 11203
rect 2329 11101 2363 11135
rect 8033 11101 8067 11135
rect 9045 11101 9079 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 12265 11101 12299 11135
rect 15393 11101 15427 11135
rect 19073 11101 19107 11135
rect 21189 11101 21223 11135
rect 21833 11101 21867 11135
rect 23581 11101 23615 11135
rect 15853 11033 15887 11067
rect 21281 11033 21315 11067
rect 23857 11033 23891 11067
rect 24685 11033 24719 11067
rect 7849 10965 7883 10999
rect 9597 10965 9631 10999
rect 12081 10965 12115 10999
rect 12725 10965 12759 10999
rect 12817 10965 12851 10999
rect 15209 10965 15243 10999
rect 18337 10965 18371 10999
rect 18429 10965 18463 10999
rect 18889 10965 18923 10999
rect 4353 10761 4387 10795
rect 10057 10761 10091 10795
rect 10149 10761 10183 10795
rect 13277 10761 13311 10795
rect 13737 10761 13771 10795
rect 16313 10761 16347 10795
rect 17601 10761 17635 10795
rect 17877 10761 17911 10795
rect 19349 10761 19383 10795
rect 24317 10761 24351 10795
rect 24685 10761 24719 10795
rect 25237 10761 25271 10795
rect 4077 10693 4111 10727
rect 5181 10693 5215 10727
rect 7021 10693 7055 10727
rect 15200 10693 15234 10727
rect 19012 10693 19046 10727
rect 20177 10693 20211 10727
rect 3801 10625 3835 10659
rect 3985 10625 4019 10659
rect 4169 10625 4203 10659
rect 4905 10625 4939 10659
rect 5053 10625 5087 10659
rect 5273 10625 5307 10659
rect 5411 10625 5445 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 7297 10625 7331 10659
rect 7573 10625 7607 10659
rect 7840 10625 7874 10659
rect 9505 10625 9539 10659
rect 9597 10625 9631 10659
rect 9781 10625 9815 10659
rect 9873 10625 9907 10659
rect 10325 10625 10359 10659
rect 10425 10625 10459 10659
rect 10609 10625 10643 10659
rect 10701 10625 10735 10659
rect 11621 10625 11655 10659
rect 11897 10625 11931 10659
rect 12153 10625 12187 10659
rect 14197 10625 14231 10659
rect 14473 10625 14507 10659
rect 14933 10625 14967 10659
rect 17325 10625 17359 10659
rect 17693 10625 17727 10659
rect 19533 10625 19567 10659
rect 24409 10625 24443 10659
rect 24501 10625 24535 10659
rect 1409 10557 1443 10591
rect 13829 10557 13863 10591
rect 13921 10557 13955 10591
rect 14381 10557 14415 10591
rect 19257 10557 19291 10591
rect 19901 10557 19935 10591
rect 25329 10557 25363 10591
rect 25421 10557 25455 10591
rect 11805 10489 11839 10523
rect 13369 10489 13403 10523
rect 24869 10489 24903 10523
rect 2053 10421 2087 10455
rect 5549 10421 5583 10455
rect 6745 10421 6779 10455
rect 8953 10421 8987 10455
rect 14197 10421 14231 10455
rect 14657 10421 14691 10455
rect 16957 10421 16991 10455
rect 17233 10421 17267 10455
rect 17417 10421 17451 10455
rect 21649 10421 21683 10455
rect 6101 10217 6135 10251
rect 6285 10217 6319 10251
rect 7941 10217 7975 10251
rect 10701 10217 10735 10251
rect 13093 10217 13127 10251
rect 13737 10217 13771 10251
rect 16865 10217 16899 10251
rect 17509 10217 17543 10251
rect 25145 10217 25179 10251
rect 6653 10149 6687 10183
rect 2513 10081 2547 10115
rect 2697 10081 2731 10115
rect 3525 10081 3559 10115
rect 4721 10081 4755 10115
rect 5641 10081 5675 10115
rect 7205 10081 7239 10115
rect 8493 10081 8527 10115
rect 9321 10081 9355 10115
rect 14841 10081 14875 10115
rect 19073 10081 19107 10115
rect 21465 10081 21499 10115
rect 21741 10081 21775 10115
rect 1501 10013 1535 10047
rect 2421 10013 2455 10047
rect 3249 10013 3283 10047
rect 3985 10013 4019 10047
rect 5365 10013 5399 10047
rect 6009 10013 6043 10047
rect 6101 10013 6135 10047
rect 6561 10013 6595 10047
rect 8309 10013 8343 10047
rect 9045 10013 9079 10047
rect 11713 10013 11747 10047
rect 13185 10013 13219 10047
rect 13369 10013 13403 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14565 10013 14599 10047
rect 14657 10013 14691 10047
rect 16313 10013 16347 10047
rect 16589 10013 16623 10047
rect 16681 10013 16715 10047
rect 16957 10013 16991 10047
rect 17049 10013 17083 10047
rect 17233 10013 17267 10047
rect 17325 10013 17359 10047
rect 23489 10013 23523 10047
rect 24869 10013 24903 10047
rect 25053 10013 25087 10047
rect 25329 10013 25363 10047
rect 25513 10013 25547 10047
rect 26525 10013 26559 10047
rect 1685 9945 1719 9979
rect 4445 9945 4479 9979
rect 5825 9945 5859 9979
rect 7021 9945 7055 9979
rect 9566 9945 9600 9979
rect 11980 9945 12014 9979
rect 15108 9945 15142 9979
rect 16497 9945 16531 9979
rect 18806 9945 18840 9979
rect 23397 9945 23431 9979
rect 2053 9877 2087 9911
rect 2881 9877 2915 9911
rect 3341 9877 3375 9911
rect 3801 9877 3835 9911
rect 4077 9877 4111 9911
rect 4537 9877 4571 9911
rect 4997 9877 5031 9911
rect 5457 9877 5491 9911
rect 6377 9877 6411 9911
rect 7113 9877 7147 9911
rect 8401 9877 8435 9911
rect 9229 9877 9263 9911
rect 14105 9877 14139 9911
rect 16221 9877 16255 9911
rect 17693 9877 17727 9911
rect 23213 9877 23247 9911
rect 24961 9877 24995 9911
rect 26341 9877 26375 9911
rect 3341 9673 3375 9707
rect 4905 9673 4939 9707
rect 7849 9673 7883 9707
rect 10885 9673 10919 9707
rect 14657 9673 14691 9707
rect 15301 9673 15335 9707
rect 15945 9673 15979 9707
rect 17693 9673 17727 9707
rect 18429 9673 18463 9707
rect 5733 9605 5767 9639
rect 8217 9605 8251 9639
rect 10241 9605 10275 9639
rect 18337 9605 18371 9639
rect 21925 9605 21959 9639
rect 24935 9605 24969 9639
rect 1869 9537 1903 9571
rect 1961 9537 1995 9571
rect 2228 9537 2262 9571
rect 3525 9537 3559 9571
rect 3792 9537 3826 9571
rect 4997 9537 5031 9571
rect 6009 9537 6043 9571
rect 6377 9537 6411 9571
rect 6633 9537 6667 9571
rect 8309 9537 8343 9571
rect 8953 9537 8987 9571
rect 9505 9537 9539 9571
rect 14105 9537 14139 9571
rect 14197 9537 14231 9571
rect 14381 9537 14415 9571
rect 14473 9537 14507 9571
rect 15485 9537 15519 9571
rect 16037 9537 16071 9571
rect 17141 9537 17175 9571
rect 17233 9537 17267 9571
rect 17417 9537 17451 9571
rect 17509 9537 17543 9571
rect 17785 9537 17819 9571
rect 21649 9537 21683 9571
rect 22017 9537 22051 9571
rect 23121 9537 23155 9571
rect 24685 9537 24719 9571
rect 24777 9537 24811 9571
rect 25053 9537 25087 9571
rect 25145 9537 25179 9571
rect 25237 9537 25271 9571
rect 25513 9537 25547 9571
rect 25605 9537 25639 9571
rect 25789 9537 25823 9571
rect 8493 9469 8527 9503
rect 10977 9469 11011 9503
rect 11069 9469 11103 9503
rect 16221 9469 16255 9503
rect 18245 9469 18279 9503
rect 21465 9469 21499 9503
rect 22753 9469 22787 9503
rect 23213 9469 23247 9503
rect 6193 9401 6227 9435
rect 10517 9401 10551 9435
rect 15577 9401 15611 9435
rect 18797 9401 18831 9435
rect 1685 9333 1719 9367
rect 7757 9333 7791 9367
rect 17969 9333 18003 9367
rect 24593 9333 24627 9367
rect 25421 9333 25455 9367
rect 25789 9333 25823 9367
rect 2973 9129 3007 9163
rect 5181 9129 5215 9163
rect 7297 9129 7331 9163
rect 13553 9129 13587 9163
rect 16957 9129 16991 9163
rect 24409 9129 24443 9163
rect 25329 9129 25363 9163
rect 2881 9061 2915 9095
rect 23489 9061 23523 9095
rect 24225 9061 24259 9095
rect 25145 9061 25179 9095
rect 3801 8993 3835 9027
rect 11161 8993 11195 9027
rect 11345 8993 11379 9027
rect 18337 8993 18371 9027
rect 21465 8993 21499 9027
rect 23213 8993 23247 9027
rect 24593 8993 24627 9027
rect 24961 8993 24995 9027
rect 1501 8925 1535 8959
rect 1768 8925 1802 8959
rect 3157 8925 3191 8959
rect 3433 8925 3467 8959
rect 5733 8925 5767 8959
rect 5917 8925 5951 8959
rect 9505 8925 9539 8959
rect 9781 8925 9815 8959
rect 13001 8925 13035 8959
rect 13369 8925 13403 8959
rect 14841 8925 14875 8959
rect 18070 8925 18104 8959
rect 23121 8925 23155 8959
rect 23581 8925 23615 8959
rect 23674 8925 23708 8959
rect 23949 8925 23983 8959
rect 24087 8925 24121 8959
rect 24685 8925 24719 8959
rect 25329 8925 25363 8959
rect 25421 8925 25455 8959
rect 25605 8925 25639 8959
rect 25881 8925 25915 8959
rect 4046 8857 4080 8891
rect 6184 8857 6218 8891
rect 10609 8857 10643 8891
rect 13185 8857 13219 8891
rect 13277 8857 13311 8891
rect 20729 8857 20763 8891
rect 21925 8857 21959 8891
rect 22293 8857 22327 8891
rect 23857 8857 23891 8891
rect 25053 8857 25087 8891
rect 3617 8789 3651 8823
rect 10701 8789 10735 8823
rect 11069 8789 11103 8823
rect 25789 8789 25823 8823
rect 8953 8585 8987 8619
rect 10517 8585 10551 8619
rect 14473 8585 14507 8619
rect 17509 8585 17543 8619
rect 17877 8585 17911 8619
rect 21557 8585 21591 8619
rect 23673 8585 23707 8619
rect 5181 8517 5215 8551
rect 9290 8517 9324 8551
rect 15301 8517 15335 8551
rect 18705 8517 18739 8551
rect 20453 8517 20487 8551
rect 20637 8517 20671 8551
rect 22477 8517 22511 8551
rect 4905 8449 4939 8483
rect 7297 8449 7331 8483
rect 8769 8449 8803 8483
rect 9045 8449 9079 8483
rect 10701 8449 10735 8483
rect 10793 8449 10827 8483
rect 10977 8449 11011 8483
rect 11069 8449 11103 8483
rect 12633 8449 12667 8483
rect 13093 8449 13127 8483
rect 13360 8449 13394 8483
rect 14565 8449 14599 8483
rect 15761 8449 15795 8483
rect 17417 8449 17451 8483
rect 19257 8449 19291 8483
rect 19717 8449 19751 8483
rect 21281 8449 21315 8483
rect 21649 8449 21683 8483
rect 22293 8449 22327 8483
rect 23305 8449 23339 8483
rect 6009 8381 6043 8415
rect 12725 8381 12759 8415
rect 12909 8381 12943 8415
rect 17325 8381 17359 8415
rect 19441 8381 19475 8415
rect 19901 8381 19935 8415
rect 20085 8381 20119 8415
rect 22017 8381 22051 8415
rect 23397 8381 23431 8415
rect 10425 8313 10459 8347
rect 15577 8313 15611 8347
rect 20269 8313 20303 8347
rect 7113 8245 7147 8279
rect 12265 8245 12299 8279
rect 20453 8245 20487 8279
rect 22753 8245 22787 8279
rect 11437 8041 11471 8075
rect 11713 8041 11747 8075
rect 13553 8041 13587 8075
rect 15945 8041 15979 8075
rect 17325 8041 17359 8075
rect 17601 8041 17635 8075
rect 20821 8041 20855 8075
rect 23765 8041 23799 8075
rect 13461 7973 13495 8007
rect 19349 7973 19383 8007
rect 9413 7905 9447 7939
rect 12081 7905 12115 7939
rect 14565 7905 14599 7939
rect 14657 7905 14691 7939
rect 16405 7905 16439 7939
rect 16497 7905 16531 7939
rect 20637 7905 20671 7939
rect 21465 7905 21499 7939
rect 21925 7905 21959 7939
rect 22109 7905 22143 7939
rect 23305 7905 23339 7939
rect 26525 7905 26559 7939
rect 6745 7837 6779 7871
rect 7012 7837 7046 7871
rect 9137 7837 9171 7871
rect 10885 7837 10919 7871
rect 11069 7837 11103 7871
rect 11253 7837 11287 7871
rect 11529 7837 11563 7871
rect 11805 7837 11839 7871
rect 13737 7837 13771 7871
rect 14473 7837 14507 7871
rect 15853 7837 15887 7871
rect 16773 7837 16807 7871
rect 17049 7837 17083 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 19717 7837 19751 7871
rect 19809 7837 19843 7871
rect 20177 7837 20211 7871
rect 20269 7837 20303 7871
rect 21281 7837 21315 7871
rect 21741 7837 21775 7871
rect 22201 7837 22235 7871
rect 23397 7837 23431 7871
rect 24501 7837 24535 7871
rect 9658 7769 9692 7803
rect 11161 7769 11195 7803
rect 12326 7769 12360 7803
rect 15025 7769 15059 7803
rect 16313 7769 16347 7803
rect 16957 7769 16991 7803
rect 22937 7769 22971 7803
rect 24777 7769 24811 7803
rect 8125 7701 8159 7735
rect 9321 7701 9355 7735
rect 10793 7701 10827 7735
rect 11989 7701 12023 7735
rect 14105 7701 14139 7735
rect 2605 7497 2639 7531
rect 5457 7497 5491 7531
rect 7297 7497 7331 7531
rect 7665 7497 7699 7531
rect 9689 7497 9723 7531
rect 10057 7497 10091 7531
rect 13185 7497 13219 7531
rect 13277 7497 13311 7531
rect 13645 7497 13679 7531
rect 13737 7497 13771 7531
rect 14381 7497 14415 7531
rect 16497 7497 16531 7531
rect 17049 7497 17083 7531
rect 17141 7497 17175 7531
rect 23121 7497 23155 7531
rect 26525 7497 26559 7531
rect 3433 7429 3467 7463
rect 4077 7429 4111 7463
rect 4169 7429 4203 7463
rect 10149 7429 10183 7463
rect 12072 7429 12106 7463
rect 15362 7429 15396 7463
rect 19901 7429 19935 7463
rect 2697 7361 2731 7395
rect 3893 7361 3927 7395
rect 4261 7361 4295 7395
rect 5273 7361 5307 7395
rect 7021 7361 7055 7395
rect 8125 7361 8159 7395
rect 8218 7361 8252 7395
rect 8401 7361 8435 7395
rect 8493 7361 8527 7395
rect 8590 7361 8624 7395
rect 14197 7361 14231 7395
rect 14841 7361 14875 7395
rect 15117 7361 15151 7395
rect 18889 7361 18923 7395
rect 18981 7361 19015 7395
rect 19441 7361 19475 7395
rect 19625 7361 19659 7395
rect 20361 7361 20395 7395
rect 20453 7361 20487 7395
rect 20913 7361 20947 7395
rect 21465 7361 21499 7395
rect 21649 7361 21683 7395
rect 22477 7361 22511 7395
rect 22661 7361 22695 7395
rect 22753 7361 22787 7395
rect 23489 7361 23523 7395
rect 23765 7361 23799 7395
rect 25053 7361 25087 7395
rect 26341 7361 26375 7395
rect 2881 7293 2915 7327
rect 3525 7293 3559 7327
rect 3709 7293 3743 7327
rect 7757 7293 7791 7327
rect 7849 7293 7883 7327
rect 10333 7293 10367 7327
rect 11805 7293 11839 7327
rect 13829 7293 13863 7327
rect 17325 7293 17359 7327
rect 18429 7293 18463 7327
rect 19809 7293 19843 7327
rect 20821 7293 20855 7327
rect 21281 7293 21315 7327
rect 22937 7293 22971 7327
rect 24685 7293 24719 7327
rect 25145 7293 25179 7327
rect 3065 7225 3099 7259
rect 21649 7225 21683 7259
rect 2237 7157 2271 7191
rect 4445 7157 4479 7191
rect 6837 7157 6871 7191
rect 8769 7157 8803 7191
rect 16681 7157 16715 7191
rect 7941 6953 7975 6987
rect 16405 6953 16439 6987
rect 19349 6953 19383 6987
rect 22477 6953 22511 6987
rect 25237 6953 25271 6987
rect 7849 6885 7883 6919
rect 8493 6817 8527 6851
rect 18245 6817 18279 6851
rect 24685 6817 24719 6851
rect 24961 6817 24995 6851
rect 25697 6817 25731 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 3433 6749 3467 6783
rect 3801 6749 3835 6783
rect 5273 6749 5307 6783
rect 5366 6749 5400 6783
rect 5641 6749 5675 6783
rect 5779 6749 5813 6783
rect 6469 6749 6503 6783
rect 6736 6749 6770 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 10057 6749 10091 6783
rect 15025 6749 15059 6783
rect 15292 6749 15326 6783
rect 18337 6749 18371 6783
rect 18521 6749 18555 6783
rect 19073 6749 19107 6783
rect 19809 6749 19843 6783
rect 19993 6749 20027 6783
rect 20269 6749 20303 6783
rect 20453 6749 20487 6783
rect 20637 6749 20671 6783
rect 21189 6749 21223 6783
rect 21281 6749 21315 6783
rect 21649 6749 21683 6783
rect 21741 6749 21775 6783
rect 22109 6749 22143 6783
rect 22201 6749 22235 6783
rect 24593 6749 24627 6783
rect 25053 6749 25087 6783
rect 25237 6749 25271 6783
rect 25513 6749 25547 6783
rect 25605 6749 25639 6783
rect 25789 6749 25823 6783
rect 2206 6681 2240 6715
rect 4046 6681 4080 6715
rect 5549 6681 5583 6715
rect 18705 6681 18739 6715
rect 22468 6681 22502 6715
rect 22845 6681 22879 6715
rect 1593 6613 1627 6647
rect 1869 6613 1903 6647
rect 3341 6613 3375 6647
rect 3617 6613 3651 6647
rect 5181 6613 5215 6647
rect 5917 6613 5951 6647
rect 9873 6613 9907 6647
rect 21005 6613 21039 6647
rect 4353 6409 4387 6443
rect 4721 6409 4755 6443
rect 4813 6409 4847 6443
rect 7757 6409 7791 6443
rect 8217 6409 8251 6443
rect 9413 6409 9447 6443
rect 10885 6409 10919 6443
rect 12909 6409 12943 6443
rect 13369 6409 13403 6443
rect 13461 6409 13495 6443
rect 19993 6409 20027 6443
rect 21189 6409 21223 6443
rect 22661 6409 22695 6443
rect 23305 6409 23339 6443
rect 23581 6409 23615 6443
rect 25437 6409 25471 6443
rect 25881 6409 25915 6443
rect 2206 6341 2240 6375
rect 3801 6341 3835 6375
rect 8309 6341 8343 6375
rect 8953 6341 8987 6375
rect 18245 6341 18279 6375
rect 21357 6341 21391 6375
rect 21557 6341 21591 6375
rect 23489 6341 23523 6375
rect 25237 6341 25271 6375
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 3893 6273 3927 6307
rect 6377 6273 6411 6307
rect 6644 6273 6678 6307
rect 9229 6273 9263 6307
rect 9505 6273 9539 6307
rect 9772 6273 9806 6307
rect 11796 6273 11830 6307
rect 18705 6273 18739 6307
rect 18797 6273 18831 6307
rect 19257 6273 19291 6307
rect 20177 6273 20211 6307
rect 20269 6273 20303 6307
rect 20729 6273 20763 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 22293 6273 22327 6307
rect 22477 6273 22511 6307
rect 22845 6273 22879 6307
rect 23121 6273 23155 6307
rect 23673 6273 23707 6307
rect 23857 6273 23891 6307
rect 24133 6273 24167 6307
rect 24225 6273 24259 6307
rect 24409 6273 24443 6307
rect 24777 6273 24811 6307
rect 25697 6273 25731 6307
rect 25973 6273 26007 6307
rect 26065 6273 26099 6307
rect 26249 6273 26283 6307
rect 4077 6205 4111 6239
rect 4997 6205 5031 6239
rect 8493 6205 8527 6239
rect 9045 6205 9079 6239
rect 11529 6205 11563 6239
rect 13645 6205 13679 6239
rect 19165 6205 19199 6239
rect 19625 6205 19659 6239
rect 20637 6205 20671 6239
rect 21097 6205 21131 6239
rect 22753 6205 22787 6239
rect 23949 6205 23983 6239
rect 24317 6205 24351 6239
rect 24869 6205 24903 6239
rect 3433 6137 3467 6171
rect 25697 6137 25731 6171
rect 1869 6069 1903 6103
rect 3341 6069 3375 6103
rect 7849 6069 7883 6103
rect 8953 6069 8987 6103
rect 13001 6069 13035 6103
rect 21373 6069 21407 6103
rect 21833 6069 21867 6103
rect 25145 6069 25179 6103
rect 25421 6069 25455 6103
rect 25605 6069 25639 6103
rect 26065 6069 26099 6103
rect 3065 5865 3099 5899
rect 6745 5865 6779 5899
rect 8217 5865 8251 5899
rect 9873 5865 9907 5899
rect 11897 5865 11931 5899
rect 19349 5865 19383 5899
rect 24041 5865 24075 5899
rect 13461 5797 13495 5831
rect 17785 5797 17819 5831
rect 1685 5729 1719 5763
rect 10517 5729 10551 5763
rect 14565 5729 14599 5763
rect 14749 5729 14783 5763
rect 16221 5729 16255 5763
rect 16313 5729 16347 5763
rect 20637 5729 20671 5763
rect 20729 5729 20763 5763
rect 24869 5729 24903 5763
rect 25053 5729 25087 5763
rect 25697 5729 25731 5763
rect 25789 5729 25823 5763
rect 1941 5661 1975 5695
rect 6929 5661 6963 5695
rect 8401 5661 8435 5695
rect 10241 5661 10275 5695
rect 12081 5661 12115 5695
rect 13645 5661 13679 5695
rect 18245 5661 18279 5695
rect 18429 5661 18463 5695
rect 18705 5661 18739 5695
rect 18889 5661 18923 5695
rect 19073 5661 19107 5695
rect 19809 5661 19843 5695
rect 19993 5661 20027 5695
rect 20177 5661 20211 5695
rect 20269 5661 20303 5695
rect 20913 5661 20947 5695
rect 21097 5661 21131 5695
rect 21557 5661 21591 5695
rect 21649 5661 21683 5695
rect 22477 5661 22511 5695
rect 22569 5661 22603 5695
rect 22661 5661 22695 5695
rect 22845 5661 22879 5695
rect 24225 5661 24259 5695
rect 24777 5661 24811 5695
rect 25605 5661 25639 5695
rect 10333 5525 10367 5559
rect 14105 5525 14139 5559
rect 14473 5525 14507 5559
rect 16405 5525 16439 5559
rect 16773 5525 16807 5559
rect 21833 5525 21867 5559
rect 22201 5525 22235 5559
rect 24409 5525 24443 5559
rect 25237 5525 25271 5559
rect 4537 5321 4571 5355
rect 5365 5321 5399 5355
rect 8309 5321 8343 5355
rect 15025 5321 15059 5355
rect 16497 5321 16531 5355
rect 16681 5321 16715 5355
rect 7941 5253 7975 5287
rect 15384 5253 15418 5287
rect 18061 5253 18095 5287
rect 19717 5253 19751 5287
rect 4445 5185 4479 5219
rect 5273 5185 5307 5219
rect 7665 5185 7699 5219
rect 7813 5185 7847 5219
rect 8033 5185 8067 5219
rect 8130 5185 8164 5219
rect 9965 5185 9999 5219
rect 13185 5185 13219 5219
rect 13369 5185 13403 5219
rect 13645 5185 13679 5219
rect 13901 5185 13935 5219
rect 16865 5185 16899 5219
rect 18245 5185 18279 5219
rect 18797 5185 18831 5219
rect 18981 5185 19015 5219
rect 19257 5185 19291 5219
rect 20269 5185 20303 5219
rect 20453 5185 20487 5219
rect 20729 5185 20763 5219
rect 4629 5117 4663 5151
rect 5457 5117 5491 5151
rect 10057 5117 10091 5151
rect 10149 5117 10183 5151
rect 15117 5117 15151 5151
rect 19165 5117 19199 5151
rect 19625 5117 19659 5151
rect 20913 5117 20947 5151
rect 21097 5117 21131 5151
rect 13553 5049 13587 5083
rect 4077 4981 4111 5015
rect 4905 4981 4939 5015
rect 9597 4981 9631 5015
rect 13001 4981 13035 5015
rect 17785 4981 17819 5015
rect 6009 4777 6043 4811
rect 6929 4777 6963 4811
rect 9413 4777 9447 4811
rect 14749 4777 14783 4811
rect 16681 4777 16715 4811
rect 10609 4709 10643 4743
rect 13921 4709 13955 4743
rect 18521 4709 18555 4743
rect 8033 4641 8067 4675
rect 10057 4641 10091 4675
rect 20729 4641 20763 4675
rect 3985 4573 4019 4607
rect 4721 4573 4755 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 5733 4573 5767 4607
rect 5825 4573 5859 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 6745 4573 6779 4607
rect 9137 4573 9171 4607
rect 9597 4573 9631 4607
rect 9781 4573 9815 4607
rect 10885 4573 10919 4607
rect 11253 4573 11287 4607
rect 12541 4573 12575 4607
rect 14105 4573 14139 4607
rect 14198 4573 14232 4607
rect 14473 4573 14507 4607
rect 14611 4573 14645 4607
rect 16819 4573 16853 4607
rect 17049 4573 17083 4607
rect 17232 4573 17266 4607
rect 17325 4573 17359 4607
rect 18981 4573 19015 4607
rect 19809 4573 19843 4607
rect 19993 4573 20027 4607
rect 20177 4573 20211 4607
rect 20269 4573 20303 4607
rect 20637 4573 20671 4607
rect 20913 4573 20947 4607
rect 21925 4573 21959 4607
rect 22201 4573 22235 4607
rect 22385 4573 22419 4607
rect 22477 4573 22511 4607
rect 23765 4573 23799 4607
rect 24593 4573 24627 4607
rect 6653 4505 6687 4539
rect 7849 4505 7883 4539
rect 10149 4505 10183 4539
rect 10977 4505 11011 4539
rect 11069 4505 11103 4539
rect 12808 4505 12842 4539
rect 14381 4505 14415 4539
rect 16957 4505 16991 4539
rect 18889 4505 18923 4539
rect 3801 4437 3835 4471
rect 4537 4437 4571 4471
rect 7481 4437 7515 4471
rect 7941 4437 7975 4471
rect 9321 4437 9355 4471
rect 10241 4437 10275 4471
rect 10701 4437 10735 4471
rect 19533 4437 19567 4471
rect 21097 4437 21131 4471
rect 21741 4437 21775 4471
rect 22569 4437 22603 4471
rect 23581 4437 23615 4471
rect 24409 4437 24443 4471
rect 5457 4233 5491 4267
rect 6837 4233 6871 4267
rect 8309 4233 8343 4267
rect 9413 4233 9447 4267
rect 13093 4233 13127 4267
rect 13461 4233 13495 4267
rect 13921 4233 13955 4267
rect 16129 4233 16163 4267
rect 17509 4233 17543 4267
rect 20085 4233 20119 4267
rect 2872 4165 2906 4199
rect 4344 4165 4378 4199
rect 9045 4165 9079 4199
rect 14289 4165 14323 4199
rect 22109 4165 22143 4199
rect 24317 4165 24351 4199
rect 2605 4097 2639 4131
rect 4077 4097 4111 4131
rect 5825 4097 5859 4131
rect 6653 4097 6687 4131
rect 7185 4097 7219 4131
rect 8953 4097 8987 4131
rect 10618 4097 10652 4131
rect 10885 4097 10919 4131
rect 11161 4097 11195 4131
rect 12633 4097 12667 4131
rect 13553 4097 13587 4131
rect 14105 4097 14139 4131
rect 14197 4097 14231 4131
rect 14473 4097 14507 4131
rect 16037 4097 16071 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 17785 4097 17819 4131
rect 17877 4097 17911 4131
rect 18061 4097 18095 4131
rect 18981 4097 19015 4131
rect 19073 4097 19107 4131
rect 19533 4097 19567 4131
rect 19717 4097 19751 4131
rect 19901 4097 19935 4131
rect 20085 4097 20119 4131
rect 20545 4097 20579 4131
rect 23857 4097 23891 4131
rect 26065 4097 26099 4131
rect 6929 4029 6963 4063
rect 8861 4029 8895 4063
rect 13645 4029 13679 4063
rect 16313 4029 16347 4063
rect 17141 4029 17175 4063
rect 17325 4029 17359 4063
rect 21833 4029 21867 4063
rect 24041 4029 24075 4063
rect 3985 3893 4019 3927
rect 5641 3893 5675 3927
rect 9505 3893 9539 3927
rect 10977 3893 11011 3927
rect 12449 3893 12483 3927
rect 15669 3893 15703 3927
rect 16681 3893 16715 3927
rect 18613 3893 18647 3927
rect 6561 3689 6595 3723
rect 8217 3689 8251 3723
rect 13553 3689 13587 3723
rect 16405 3689 16439 3723
rect 17877 3689 17911 3723
rect 24961 3689 24995 3723
rect 10609 3621 10643 3655
rect 18705 3621 18739 3655
rect 9229 3553 9263 3587
rect 12173 3553 12207 3587
rect 14565 3553 14599 3587
rect 14749 3553 14783 3587
rect 18153 3553 18187 3587
rect 21097 3553 21131 3587
rect 21373 3553 21407 3587
rect 21741 3553 21775 3587
rect 23489 3553 23523 3587
rect 4721 3485 4755 3519
rect 5181 3485 5215 3519
rect 6837 3485 6871 3519
rect 8953 3485 8987 3519
rect 9485 3485 9519 3519
rect 11897 3485 11931 3519
rect 12440 3485 12474 3519
rect 14473 3485 14507 3519
rect 15025 3485 15059 3519
rect 16497 3485 16531 3519
rect 18981 3485 19015 3519
rect 21005 3485 21039 3519
rect 21465 3485 21499 3519
rect 24593 3485 24627 3519
rect 24869 3485 24903 3519
rect 5448 3417 5482 3451
rect 7104 3417 7138 3451
rect 15292 3417 15326 3451
rect 16742 3417 16776 3451
rect 4537 3349 4571 3383
rect 9137 3349 9171 3383
rect 12081 3349 12115 3383
rect 14105 3349 14139 3383
rect 18245 3349 18279 3383
rect 18337 3349 18371 3383
rect 18797 3349 18831 3383
rect 24501 3349 24535 3383
rect 5457 3145 5491 3179
rect 5825 3145 5859 3179
rect 6377 3145 6411 3179
rect 6745 3145 6779 3179
rect 7205 3145 7239 3179
rect 7481 3145 7515 3179
rect 7849 3145 7883 3179
rect 10609 3145 10643 3179
rect 13277 3145 13311 3179
rect 13369 3145 13403 3179
rect 13737 3145 13771 3179
rect 15393 3145 15427 3179
rect 16313 3145 16347 3179
rect 17049 3145 17083 3179
rect 22569 3145 22603 3179
rect 24869 3145 24903 3179
rect 9474 3077 9508 3111
rect 18184 3077 18218 3111
rect 23397 3077 23431 3111
rect 3985 3009 4019 3043
rect 4252 3009 4286 3043
rect 5917 3009 5951 3043
rect 6837 3009 6871 3043
rect 7389 3009 7423 3043
rect 7941 3009 7975 3043
rect 9229 3009 9263 3043
rect 11897 3009 11931 3043
rect 12164 3009 12198 3043
rect 13829 3009 13863 3043
rect 15577 3009 15611 3043
rect 16129 3009 16163 3043
rect 22477 3009 22511 3043
rect 6101 2941 6135 2975
rect 7021 2941 7055 2975
rect 8125 2941 8159 2975
rect 14013 2941 14047 2975
rect 18429 2941 18463 2975
rect 23121 2941 23155 2975
rect 5365 2805 5399 2839
rect 6009 2601 6043 2635
rect 16221 2533 16255 2567
rect 9229 2465 9263 2499
rect 13277 2465 13311 2499
rect 6929 2397 6963 2431
rect 8217 2397 8251 2431
rect 8769 2397 8803 2431
rect 8953 2397 8987 2431
rect 12357 2397 12391 2431
rect 12909 2397 12943 2431
rect 13001 2397 13035 2431
rect 17233 2397 17267 2431
rect 6101 2329 6135 2363
rect 6377 2329 6411 2363
rect 16405 2329 16439 2363
rect 16681 2329 16715 2363
<< metal1 >>
rect 1104 27770 26864 27792
rect 1104 27718 2918 27770
rect 2970 27718 2982 27770
rect 3034 27718 3046 27770
rect 3098 27718 3110 27770
rect 3162 27718 3174 27770
rect 3226 27718 3238 27770
rect 3290 27718 6918 27770
rect 6970 27718 6982 27770
rect 7034 27718 7046 27770
rect 7098 27718 7110 27770
rect 7162 27718 7174 27770
rect 7226 27718 7238 27770
rect 7290 27718 10918 27770
rect 10970 27718 10982 27770
rect 11034 27718 11046 27770
rect 11098 27718 11110 27770
rect 11162 27718 11174 27770
rect 11226 27718 11238 27770
rect 11290 27718 14918 27770
rect 14970 27718 14982 27770
rect 15034 27718 15046 27770
rect 15098 27718 15110 27770
rect 15162 27718 15174 27770
rect 15226 27718 15238 27770
rect 15290 27718 18918 27770
rect 18970 27718 18982 27770
rect 19034 27718 19046 27770
rect 19098 27718 19110 27770
rect 19162 27718 19174 27770
rect 19226 27718 19238 27770
rect 19290 27718 22918 27770
rect 22970 27718 22982 27770
rect 23034 27718 23046 27770
rect 23098 27718 23110 27770
rect 23162 27718 23174 27770
rect 23226 27718 23238 27770
rect 23290 27718 26864 27770
rect 1104 27696 26864 27718
rect 9766 27548 9772 27600
rect 9824 27548 9830 27600
rect 10318 27548 10324 27600
rect 10376 27588 10382 27600
rect 10413 27591 10471 27597
rect 10413 27588 10425 27591
rect 10376 27560 10425 27588
rect 10376 27548 10382 27560
rect 10413 27557 10425 27560
rect 10459 27557 10471 27591
rect 10413 27551 10471 27557
rect 10778 27548 10784 27600
rect 10836 27588 10842 27600
rect 11057 27591 11115 27597
rect 11057 27588 11069 27591
rect 10836 27560 11069 27588
rect 10836 27548 10842 27560
rect 11057 27557 11069 27560
rect 11103 27557 11115 27591
rect 11057 27551 11115 27557
rect 11698 27548 11704 27600
rect 11756 27548 11762 27600
rect 12342 27548 12348 27600
rect 12400 27548 12406 27600
rect 14274 27548 14280 27600
rect 14332 27548 14338 27600
rect 17402 27548 17408 27600
rect 17460 27588 17466 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 17460 27560 17509 27588
rect 17460 27548 17466 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 17497 27551 17555 27557
rect 20070 27548 20076 27600
rect 20128 27548 20134 27600
rect 20622 27480 20628 27532
rect 20680 27520 20686 27532
rect 20717 27523 20775 27529
rect 20717 27520 20729 27523
rect 20680 27492 20729 27520
rect 20680 27480 20686 27492
rect 20717 27489 20729 27492
rect 20763 27489 20775 27523
rect 20717 27483 20775 27489
rect 9766 27412 9772 27464
rect 9824 27452 9830 27464
rect 9953 27455 10011 27461
rect 9953 27452 9965 27455
rect 9824 27424 9965 27452
rect 9824 27412 9830 27424
rect 9953 27421 9965 27424
rect 9999 27421 10011 27455
rect 9953 27415 10011 27421
rect 10594 27412 10600 27464
rect 10652 27412 10658 27464
rect 11241 27455 11299 27461
rect 11241 27421 11253 27455
rect 11287 27452 11299 27455
rect 11514 27452 11520 27464
rect 11287 27424 11520 27452
rect 11287 27421 11299 27424
rect 11241 27415 11299 27421
rect 11514 27412 11520 27424
rect 11572 27412 11578 27464
rect 11885 27455 11943 27461
rect 11885 27421 11897 27455
rect 11931 27421 11943 27455
rect 11885 27415 11943 27421
rect 11422 27344 11428 27396
rect 11480 27384 11486 27396
rect 11900 27384 11928 27415
rect 12158 27412 12164 27464
rect 12216 27452 12222 27464
rect 12529 27455 12587 27461
rect 12529 27452 12541 27455
rect 12216 27424 12541 27452
rect 12216 27412 12222 27424
rect 12529 27421 12541 27424
rect 12575 27421 12587 27455
rect 12529 27415 12587 27421
rect 14458 27412 14464 27464
rect 14516 27412 14522 27464
rect 17678 27412 17684 27464
rect 17736 27412 17742 27464
rect 19426 27412 19432 27464
rect 19484 27412 19490 27464
rect 19518 27412 19524 27464
rect 19576 27452 19582 27464
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 19576 27424 19625 27452
rect 19576 27412 19582 27424
rect 19613 27421 19625 27424
rect 19659 27421 19671 27455
rect 19613 27415 19671 27421
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27452 19763 27455
rect 20070 27452 20076 27464
rect 19751 27424 20076 27452
rect 19751 27421 19763 27424
rect 19705 27415 19763 27421
rect 20070 27412 20076 27424
rect 20128 27412 20134 27464
rect 20257 27455 20315 27461
rect 20257 27421 20269 27455
rect 20303 27452 20315 27455
rect 20530 27452 20536 27464
rect 20303 27424 20536 27452
rect 20303 27421 20315 27424
rect 20257 27415 20315 27421
rect 20530 27412 20536 27424
rect 20588 27412 20594 27464
rect 21361 27455 21419 27461
rect 21361 27421 21373 27455
rect 21407 27452 21419 27455
rect 21453 27455 21511 27461
rect 21453 27452 21465 27455
rect 21407 27424 21465 27452
rect 21407 27421 21419 27424
rect 21361 27415 21419 27421
rect 21453 27421 21465 27424
rect 21499 27421 21511 27455
rect 21453 27415 21511 27421
rect 11480 27356 11928 27384
rect 11480 27344 11486 27356
rect 18690 27276 18696 27328
rect 18748 27316 18754 27328
rect 19245 27319 19303 27325
rect 19245 27316 19257 27319
rect 18748 27288 19257 27316
rect 18748 27276 18754 27288
rect 19245 27285 19257 27288
rect 19291 27285 19303 27319
rect 19245 27279 19303 27285
rect 21082 27276 21088 27328
rect 21140 27316 21146 27328
rect 21637 27319 21695 27325
rect 21637 27316 21649 27319
rect 21140 27288 21649 27316
rect 21140 27276 21146 27288
rect 21637 27285 21649 27288
rect 21683 27285 21695 27319
rect 21637 27279 21695 27285
rect 1104 27226 26864 27248
rect 1104 27174 3658 27226
rect 3710 27174 3722 27226
rect 3774 27174 3786 27226
rect 3838 27174 3850 27226
rect 3902 27174 3914 27226
rect 3966 27174 3978 27226
rect 4030 27174 7658 27226
rect 7710 27174 7722 27226
rect 7774 27174 7786 27226
rect 7838 27174 7850 27226
rect 7902 27174 7914 27226
rect 7966 27174 7978 27226
rect 8030 27174 11658 27226
rect 11710 27174 11722 27226
rect 11774 27174 11786 27226
rect 11838 27174 11850 27226
rect 11902 27174 11914 27226
rect 11966 27174 11978 27226
rect 12030 27174 15658 27226
rect 15710 27174 15722 27226
rect 15774 27174 15786 27226
rect 15838 27174 15850 27226
rect 15902 27174 15914 27226
rect 15966 27174 15978 27226
rect 16030 27174 19658 27226
rect 19710 27174 19722 27226
rect 19774 27174 19786 27226
rect 19838 27174 19850 27226
rect 19902 27174 19914 27226
rect 19966 27174 19978 27226
rect 20030 27174 23658 27226
rect 23710 27174 23722 27226
rect 23774 27174 23786 27226
rect 23838 27174 23850 27226
rect 23902 27174 23914 27226
rect 23966 27174 23978 27226
rect 24030 27174 26864 27226
rect 1104 27152 26864 27174
rect 7929 27115 7987 27121
rect 7929 27081 7941 27115
rect 7975 27081 7987 27115
rect 7929 27075 7987 27081
rect 4982 26936 4988 26988
rect 5040 26936 5046 26988
rect 7837 26979 7895 26985
rect 7837 26945 7849 26979
rect 7883 26976 7895 26979
rect 7944 26976 7972 27075
rect 9766 27072 9772 27124
rect 9824 27112 9830 27124
rect 9824 27084 11008 27112
rect 9824 27072 9830 27084
rect 10778 27044 10784 27056
rect 10428 27016 10784 27044
rect 7883 26948 7972 26976
rect 8297 26979 8355 26985
rect 7883 26945 7895 26948
rect 7837 26939 7895 26945
rect 8297 26945 8309 26979
rect 8343 26976 8355 26979
rect 8754 26976 8760 26988
rect 8343 26948 8760 26976
rect 8343 26945 8355 26948
rect 8297 26939 8355 26945
rect 8754 26936 8760 26948
rect 8812 26936 8818 26988
rect 9769 26979 9827 26985
rect 9769 26945 9781 26979
rect 9815 26976 9827 26979
rect 9953 26979 10011 26985
rect 9815 26948 9904 26976
rect 9815 26945 9827 26948
rect 9769 26939 9827 26945
rect 8386 26868 8392 26920
rect 8444 26868 8450 26920
rect 8570 26868 8576 26920
rect 8628 26868 8634 26920
rect 9306 26868 9312 26920
rect 9364 26908 9370 26920
rect 9493 26911 9551 26917
rect 9493 26908 9505 26911
rect 9364 26880 9505 26908
rect 9364 26868 9370 26880
rect 9493 26877 9505 26880
rect 9539 26877 9551 26911
rect 9493 26871 9551 26877
rect 9674 26800 9680 26852
rect 9732 26840 9738 26852
rect 9876 26840 9904 26948
rect 9953 26945 9965 26979
rect 9999 26976 10011 26979
rect 10045 26979 10103 26985
rect 10045 26976 10057 26979
rect 9999 26948 10057 26976
rect 9999 26945 10011 26948
rect 9953 26939 10011 26945
rect 10045 26945 10057 26948
rect 10091 26945 10103 26979
rect 10045 26939 10103 26945
rect 10226 26936 10232 26988
rect 10284 26936 10290 26988
rect 10428 26985 10456 27016
rect 10778 27004 10784 27016
rect 10836 27004 10842 27056
rect 10980 27053 11008 27084
rect 11054 27072 11060 27124
rect 11112 27112 11118 27124
rect 19426 27112 19432 27124
rect 11112 27084 19432 27112
rect 11112 27072 11118 27084
rect 10965 27047 11023 27053
rect 10965 27013 10977 27047
rect 11011 27013 11023 27047
rect 10965 27007 11023 27013
rect 12526 27004 12532 27056
rect 12584 27044 12590 27056
rect 13725 27047 13783 27053
rect 13725 27044 13737 27047
rect 12584 27016 13737 27044
rect 12584 27004 12590 27016
rect 13725 27013 13737 27016
rect 13771 27013 13783 27047
rect 14461 27047 14519 27053
rect 14461 27044 14473 27047
rect 13725 27007 13783 27013
rect 13924 27016 14473 27044
rect 10321 26979 10379 26985
rect 10321 26945 10333 26979
rect 10367 26945 10379 26979
rect 10321 26939 10379 26945
rect 10413 26979 10471 26985
rect 10413 26945 10425 26979
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 10336 26908 10364 26939
rect 10686 26936 10692 26988
rect 10744 26936 10750 26988
rect 10870 26936 10876 26988
rect 10928 26936 10934 26988
rect 11057 26979 11115 26985
rect 11057 26945 11069 26979
rect 11103 26976 11115 26979
rect 11103 26948 12020 26976
rect 11103 26945 11115 26948
rect 11057 26939 11115 26945
rect 10594 26908 10600 26920
rect 10336 26880 10600 26908
rect 10594 26868 10600 26880
rect 10652 26908 10658 26920
rect 11882 26908 11888 26920
rect 10652 26880 11888 26908
rect 10652 26868 10658 26880
rect 11882 26868 11888 26880
rect 11940 26868 11946 26920
rect 11992 26908 12020 26948
rect 12986 26936 12992 26988
rect 13044 26936 13050 26988
rect 13538 26936 13544 26988
rect 13596 26936 13602 26988
rect 13924 26985 13952 27016
rect 14461 27013 14473 27016
rect 14507 27013 14519 27047
rect 14461 27007 14519 27013
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26945 13691 26979
rect 13633 26939 13691 26945
rect 13909 26979 13967 26985
rect 13909 26945 13921 26979
rect 13955 26945 13967 26979
rect 13909 26939 13967 26945
rect 14277 26979 14335 26985
rect 14277 26945 14289 26979
rect 14323 26976 14335 26979
rect 14568 26976 14596 27084
rect 14844 27016 16344 27044
rect 14844 26988 14872 27016
rect 14323 26948 14596 26976
rect 14737 26979 14795 26985
rect 14323 26945 14335 26948
rect 14277 26939 14335 26945
rect 14737 26945 14749 26979
rect 14783 26976 14795 26979
rect 14826 26976 14832 26988
rect 14783 26948 14832 26976
rect 14783 26945 14795 26948
rect 14737 26939 14795 26945
rect 13556 26908 13584 26936
rect 11992 26880 13584 26908
rect 9732 26812 10732 26840
rect 9732 26800 9738 26812
rect 4798 26732 4804 26784
rect 4856 26732 4862 26784
rect 7650 26732 7656 26784
rect 7708 26732 7714 26784
rect 9214 26732 9220 26784
rect 9272 26772 9278 26784
rect 9585 26775 9643 26781
rect 9585 26772 9597 26775
rect 9272 26744 9597 26772
rect 9272 26732 9278 26744
rect 9585 26741 9597 26744
rect 9631 26741 9643 26775
rect 9585 26735 9643 26741
rect 10502 26732 10508 26784
rect 10560 26772 10566 26784
rect 10597 26775 10655 26781
rect 10597 26772 10609 26775
rect 10560 26744 10609 26772
rect 10560 26732 10566 26744
rect 10597 26741 10609 26744
rect 10643 26741 10655 26775
rect 10704 26772 10732 26812
rect 10778 26800 10784 26852
rect 10836 26840 10842 26852
rect 11992 26840 12020 26880
rect 10836 26812 12020 26840
rect 13648 26840 13676 26939
rect 14826 26936 14832 26948
rect 14884 26936 14890 26988
rect 16316 26985 16344 27016
rect 17144 26985 17172 27084
rect 19426 27072 19432 27084
rect 19484 27112 19490 27124
rect 20898 27112 20904 27124
rect 19484 27084 20904 27112
rect 19484 27072 19490 27084
rect 20898 27072 20904 27084
rect 20956 27072 20962 27124
rect 19518 27044 19524 27056
rect 17236 27016 19524 27044
rect 17236 26988 17264 27016
rect 19518 27004 19524 27016
rect 19576 27044 19582 27056
rect 20346 27044 20352 27056
rect 19576 27016 20352 27044
rect 19576 27004 19582 27016
rect 20346 27004 20352 27016
rect 20404 27004 20410 27056
rect 15105 26979 15163 26985
rect 15105 26945 15117 26979
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 16301 26979 16359 26985
rect 16301 26945 16313 26979
rect 16347 26945 16359 26979
rect 16301 26939 16359 26945
rect 17097 26979 17172 26985
rect 17097 26945 17109 26979
rect 17143 26948 17172 26979
rect 17143 26945 17155 26948
rect 17097 26939 17155 26945
rect 13814 26868 13820 26920
rect 13872 26908 13878 26920
rect 14001 26911 14059 26917
rect 14001 26908 14013 26911
rect 13872 26880 14013 26908
rect 13872 26868 13878 26880
rect 14001 26877 14013 26880
rect 14047 26877 14059 26911
rect 15120 26908 15148 26939
rect 17218 26936 17224 26988
rect 17276 26936 17282 26988
rect 17313 26979 17371 26985
rect 17313 26945 17325 26979
rect 17359 26976 17371 26979
rect 17586 26976 17592 26988
rect 17359 26948 17592 26976
rect 17359 26945 17371 26948
rect 17313 26939 17371 26945
rect 17586 26936 17592 26948
rect 17644 26976 17650 26988
rect 17773 26979 17831 26985
rect 17773 26976 17785 26979
rect 17644 26948 17785 26976
rect 17644 26936 17650 26948
rect 17773 26945 17785 26948
rect 17819 26945 17831 26979
rect 17773 26939 17831 26945
rect 18598 26936 18604 26988
rect 18656 26976 18662 26988
rect 19041 26979 19099 26985
rect 19041 26976 19053 26979
rect 18656 26948 19053 26976
rect 18656 26936 18662 26948
rect 19041 26945 19053 26948
rect 19087 26945 19099 26979
rect 19041 26939 19099 26945
rect 20257 26979 20315 26985
rect 20257 26945 20269 26979
rect 20303 26976 20315 26979
rect 20806 26976 20812 26988
rect 20303 26948 20812 26976
rect 20303 26945 20315 26948
rect 20257 26939 20315 26945
rect 20806 26936 20812 26948
rect 20864 26936 20870 26988
rect 16574 26908 16580 26920
rect 15120 26880 16580 26908
rect 14001 26871 14059 26877
rect 16574 26868 16580 26880
rect 16632 26868 16638 26920
rect 17402 26868 17408 26920
rect 17460 26908 17466 26920
rect 17865 26911 17923 26917
rect 17865 26908 17877 26911
rect 17460 26880 17877 26908
rect 17460 26868 17466 26880
rect 17865 26877 17877 26880
rect 17911 26877 17923 26911
rect 17865 26871 17923 26877
rect 17957 26911 18015 26917
rect 17957 26877 17969 26911
rect 18003 26877 18015 26911
rect 17957 26871 18015 26877
rect 14458 26840 14464 26852
rect 13648 26812 14464 26840
rect 10836 26800 10842 26812
rect 14458 26800 14464 26812
rect 14516 26800 14522 26852
rect 16853 26843 16911 26849
rect 14568 26812 16620 26840
rect 10962 26772 10968 26784
rect 10704 26744 10968 26772
rect 10597 26735 10655 26741
rect 10962 26732 10968 26744
rect 11020 26732 11026 26784
rect 11241 26775 11299 26781
rect 11241 26741 11253 26775
rect 11287 26772 11299 26775
rect 11330 26772 11336 26784
rect 11287 26744 11336 26772
rect 11287 26741 11299 26744
rect 11241 26735 11299 26741
rect 11330 26732 11336 26744
rect 11388 26732 11394 26784
rect 12710 26732 12716 26784
rect 12768 26772 12774 26784
rect 12805 26775 12863 26781
rect 12805 26772 12817 26775
rect 12768 26744 12817 26772
rect 12768 26732 12774 26744
rect 12805 26741 12817 26744
rect 12851 26741 12863 26775
rect 12805 26735 12863 26741
rect 13354 26732 13360 26784
rect 13412 26732 13418 26784
rect 13906 26732 13912 26784
rect 13964 26772 13970 26784
rect 14093 26775 14151 26781
rect 14093 26772 14105 26775
rect 13964 26744 14105 26772
rect 13964 26732 13970 26744
rect 14093 26741 14105 26744
rect 14139 26772 14151 26775
rect 14568 26772 14596 26812
rect 14139 26744 14596 26772
rect 14139 26741 14151 26744
rect 14093 26735 14151 26741
rect 14642 26732 14648 26784
rect 14700 26732 14706 26784
rect 14734 26732 14740 26784
rect 14792 26772 14798 26784
rect 14921 26775 14979 26781
rect 14921 26772 14933 26775
rect 14792 26744 14933 26772
rect 14792 26732 14798 26744
rect 14921 26741 14933 26744
rect 14967 26741 14979 26775
rect 14921 26735 14979 26741
rect 16393 26775 16451 26781
rect 16393 26741 16405 26775
rect 16439 26772 16451 26775
rect 16482 26772 16488 26784
rect 16439 26744 16488 26772
rect 16439 26741 16451 26744
rect 16393 26735 16451 26741
rect 16482 26732 16488 26744
rect 16540 26732 16546 26784
rect 16592 26772 16620 26812
rect 16853 26809 16865 26843
rect 16899 26840 16911 26843
rect 17494 26840 17500 26852
rect 16899 26812 17500 26840
rect 16899 26809 16911 26812
rect 16853 26803 16911 26809
rect 17494 26800 17500 26812
rect 17552 26800 17558 26852
rect 17972 26840 18000 26871
rect 18782 26868 18788 26920
rect 18840 26868 18846 26920
rect 17880 26812 18000 26840
rect 17880 26784 17908 26812
rect 17218 26772 17224 26784
rect 16592 26744 17224 26772
rect 17218 26732 17224 26744
rect 17276 26732 17282 26784
rect 17402 26732 17408 26784
rect 17460 26732 17466 26784
rect 17862 26732 17868 26784
rect 17920 26732 17926 26784
rect 20070 26732 20076 26784
rect 20128 26772 20134 26784
rect 20165 26775 20223 26781
rect 20165 26772 20177 26775
rect 20128 26744 20177 26772
rect 20128 26732 20134 26744
rect 20165 26741 20177 26744
rect 20211 26741 20223 26775
rect 20165 26735 20223 26741
rect 20254 26732 20260 26784
rect 20312 26772 20318 26784
rect 20349 26775 20407 26781
rect 20349 26772 20361 26775
rect 20312 26744 20361 26772
rect 20312 26732 20318 26744
rect 20349 26741 20361 26744
rect 20395 26741 20407 26775
rect 20349 26735 20407 26741
rect 1104 26682 26864 26704
rect 1104 26630 2918 26682
rect 2970 26630 2982 26682
rect 3034 26630 3046 26682
rect 3098 26630 3110 26682
rect 3162 26630 3174 26682
rect 3226 26630 3238 26682
rect 3290 26630 6918 26682
rect 6970 26630 6982 26682
rect 7034 26630 7046 26682
rect 7098 26630 7110 26682
rect 7162 26630 7174 26682
rect 7226 26630 7238 26682
rect 7290 26630 10918 26682
rect 10970 26630 10982 26682
rect 11034 26630 11046 26682
rect 11098 26630 11110 26682
rect 11162 26630 11174 26682
rect 11226 26630 11238 26682
rect 11290 26630 14918 26682
rect 14970 26630 14982 26682
rect 15034 26630 15046 26682
rect 15098 26630 15110 26682
rect 15162 26630 15174 26682
rect 15226 26630 15238 26682
rect 15290 26630 18918 26682
rect 18970 26630 18982 26682
rect 19034 26630 19046 26682
rect 19098 26630 19110 26682
rect 19162 26630 19174 26682
rect 19226 26630 19238 26682
rect 19290 26630 22918 26682
rect 22970 26630 22982 26682
rect 23034 26630 23046 26682
rect 23098 26630 23110 26682
rect 23162 26630 23174 26682
rect 23226 26630 23238 26682
rect 23290 26630 26864 26682
rect 1104 26608 26864 26630
rect 5074 26528 5080 26580
rect 5132 26568 5138 26580
rect 5813 26571 5871 26577
rect 5813 26568 5825 26571
rect 5132 26540 5825 26568
rect 5132 26528 5138 26540
rect 5813 26537 5825 26540
rect 5859 26537 5871 26571
rect 5813 26531 5871 26537
rect 7392 26540 8340 26568
rect 7392 26500 7420 26540
rect 7300 26472 7420 26500
rect 8312 26500 8340 26540
rect 8754 26528 8760 26580
rect 8812 26568 8818 26580
rect 9030 26568 9036 26580
rect 8812 26540 9036 26568
rect 8812 26528 8818 26540
rect 9030 26528 9036 26540
rect 9088 26528 9094 26580
rect 11882 26528 11888 26580
rect 11940 26528 11946 26580
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 16724 26540 19288 26568
rect 16724 26528 16730 26540
rect 8941 26503 8999 26509
rect 8941 26500 8953 26503
rect 8312 26472 8953 26500
rect 5442 26392 5448 26444
rect 5500 26432 5506 26444
rect 7006 26432 7012 26444
rect 5500 26404 7012 26432
rect 5500 26392 5506 26404
rect 7006 26392 7012 26404
rect 7064 26432 7070 26444
rect 7190 26432 7196 26444
rect 7064 26404 7196 26432
rect 7064 26392 7070 26404
rect 7190 26392 7196 26404
rect 7248 26392 7254 26444
rect 4062 26324 4068 26376
rect 4120 26324 4126 26376
rect 4430 26364 4436 26376
rect 4391 26336 4436 26364
rect 4430 26324 4436 26336
rect 4488 26364 4494 26376
rect 5460 26364 5488 26392
rect 7300 26373 7328 26472
rect 8941 26469 8953 26472
rect 8987 26469 8999 26503
rect 8941 26463 8999 26469
rect 17586 26460 17592 26512
rect 17644 26460 17650 26512
rect 7374 26392 7380 26444
rect 7432 26392 7438 26444
rect 8570 26392 8576 26444
rect 8628 26432 8634 26444
rect 9493 26435 9551 26441
rect 9493 26432 9505 26435
rect 8628 26404 9505 26432
rect 8628 26392 8634 26404
rect 9493 26401 9505 26404
rect 9539 26401 9551 26435
rect 9493 26395 9551 26401
rect 10137 26435 10195 26441
rect 10137 26401 10149 26435
rect 10183 26432 10195 26435
rect 10410 26432 10416 26444
rect 10183 26404 10416 26432
rect 10183 26401 10195 26404
rect 10137 26395 10195 26401
rect 10410 26392 10416 26404
rect 10468 26392 10474 26444
rect 17497 26435 17555 26441
rect 15672 26404 17264 26432
rect 7650 26373 7656 26376
rect 4488 26336 5488 26364
rect 7285 26367 7343 26373
rect 4488 26324 4494 26336
rect 7285 26333 7297 26367
rect 7331 26333 7343 26367
rect 7285 26327 7343 26333
rect 7644 26327 7656 26373
rect 7708 26364 7714 26376
rect 12161 26367 12219 26373
rect 7708 26336 7744 26364
rect 7650 26324 7656 26327
rect 7708 26324 7714 26336
rect 12161 26333 12173 26367
rect 12207 26364 12219 26367
rect 12250 26364 12256 26376
rect 12207 26336 12256 26364
rect 12207 26333 12219 26336
rect 12161 26327 12219 26333
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 12434 26324 12440 26376
rect 12492 26324 12498 26376
rect 12710 26373 12716 26376
rect 12704 26364 12716 26373
rect 12671 26336 12716 26364
rect 12704 26327 12716 26336
rect 12710 26324 12716 26327
rect 12768 26324 12774 26376
rect 14090 26324 14096 26376
rect 14148 26364 14154 26376
rect 14277 26367 14335 26373
rect 14277 26364 14289 26367
rect 14148 26336 14289 26364
rect 14148 26324 14154 26336
rect 14277 26333 14289 26336
rect 14323 26364 14335 26367
rect 15672 26364 15700 26404
rect 14323 26336 15700 26364
rect 15749 26367 15807 26373
rect 14323 26333 14335 26336
rect 14277 26327 14335 26333
rect 15749 26333 15761 26367
rect 15795 26333 15807 26367
rect 17236 26364 17264 26404
rect 17497 26401 17509 26435
rect 17543 26432 17555 26435
rect 17678 26432 17684 26444
rect 17543 26404 17684 26432
rect 17543 26401 17555 26404
rect 17497 26395 17555 26401
rect 17678 26392 17684 26404
rect 17736 26392 17742 26444
rect 19260 26441 19288 26540
rect 19245 26435 19303 26441
rect 19245 26401 19257 26435
rect 19291 26401 19303 26435
rect 19245 26395 19303 26401
rect 20530 26392 20536 26444
rect 20588 26432 20594 26444
rect 20993 26435 21051 26441
rect 20993 26432 21005 26435
rect 20588 26404 21005 26432
rect 20588 26392 20594 26404
rect 20993 26401 21005 26404
rect 21039 26401 21051 26435
rect 20993 26395 21051 26401
rect 18874 26364 18880 26376
rect 17236 26336 18880 26364
rect 15749 26327 15807 26333
rect 4700 26299 4758 26305
rect 4700 26265 4712 26299
rect 4746 26296 4758 26299
rect 4798 26296 4804 26308
rect 4746 26268 4804 26296
rect 4746 26265 4758 26268
rect 4700 26259 4758 26265
rect 4798 26256 4804 26268
rect 4856 26256 4862 26308
rect 10413 26299 10471 26305
rect 10413 26265 10425 26299
rect 10459 26296 10471 26299
rect 10502 26296 10508 26308
rect 10459 26268 10508 26296
rect 10459 26265 10471 26268
rect 10413 26259 10471 26265
rect 10502 26256 10508 26268
rect 10560 26256 10566 26308
rect 12069 26299 12127 26305
rect 12069 26296 12081 26299
rect 11638 26268 12081 26296
rect 12069 26265 12081 26268
rect 12115 26265 12127 26299
rect 12069 26259 12127 26265
rect 14544 26299 14602 26305
rect 14544 26265 14556 26299
rect 14590 26296 14602 26299
rect 14734 26296 14740 26308
rect 14590 26268 14740 26296
rect 14590 26265 14602 26268
rect 14544 26259 14602 26265
rect 14734 26256 14740 26268
rect 14792 26256 14798 26308
rect 15562 26256 15568 26308
rect 15620 26296 15626 26308
rect 15764 26296 15792 26327
rect 18874 26324 18880 26336
rect 18932 26364 18938 26376
rect 18969 26367 19027 26373
rect 18969 26364 18981 26367
rect 18932 26336 18981 26364
rect 18932 26324 18938 26336
rect 18969 26333 18981 26336
rect 19015 26333 19027 26367
rect 18969 26327 19027 26333
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 21085 26367 21143 26373
rect 21085 26364 21097 26367
rect 20956 26336 21097 26364
rect 20956 26324 20962 26336
rect 21085 26333 21097 26336
rect 21131 26333 21143 26367
rect 21085 26327 21143 26333
rect 21266 26324 21272 26376
rect 21324 26324 21330 26376
rect 22094 26324 22100 26376
rect 22152 26364 22158 26376
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 22152 26336 23213 26364
rect 22152 26324 22158 26336
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 15620 26268 15792 26296
rect 16025 26299 16083 26305
rect 15620 26256 15626 26268
rect 16025 26265 16037 26299
rect 16071 26296 16083 26299
rect 16071 26268 16436 26296
rect 16071 26265 16083 26268
rect 16025 26259 16083 26265
rect 3510 26188 3516 26240
rect 3568 26228 3574 26240
rect 3881 26231 3939 26237
rect 3881 26228 3893 26231
rect 3568 26200 3893 26228
rect 3568 26188 3574 26200
rect 3881 26197 3893 26200
rect 3927 26197 3939 26231
rect 3881 26191 3939 26197
rect 7098 26188 7104 26240
rect 7156 26188 7162 26240
rect 9306 26188 9312 26240
rect 9364 26188 9370 26240
rect 9398 26188 9404 26240
rect 9456 26188 9462 26240
rect 13814 26188 13820 26240
rect 13872 26188 13878 26240
rect 15657 26231 15715 26237
rect 15657 26197 15669 26231
rect 15703 26228 15715 26231
rect 16114 26228 16120 26240
rect 15703 26200 16120 26228
rect 15703 26197 15715 26200
rect 15657 26191 15715 26197
rect 16114 26188 16120 26200
rect 16172 26188 16178 26240
rect 16408 26228 16436 26268
rect 16482 26256 16488 26308
rect 16540 26256 16546 26308
rect 17328 26268 17908 26296
rect 17328 26228 17356 26268
rect 16408 26200 17356 26228
rect 17880 26228 17908 26268
rect 17954 26256 17960 26308
rect 18012 26296 18018 26308
rect 18702 26299 18760 26305
rect 18702 26296 18714 26299
rect 18012 26268 18714 26296
rect 18012 26256 18018 26268
rect 18702 26265 18714 26268
rect 18748 26265 18760 26299
rect 18702 26259 18760 26265
rect 19518 26256 19524 26308
rect 19576 26256 19582 26308
rect 20254 26256 20260 26308
rect 20312 26256 20318 26308
rect 23293 26299 23351 26305
rect 23293 26265 23305 26299
rect 23339 26296 23351 26299
rect 23474 26296 23480 26308
rect 23339 26268 23480 26296
rect 23339 26265 23351 26268
rect 23293 26259 23351 26265
rect 23474 26256 23480 26268
rect 23532 26256 23538 26308
rect 18046 26228 18052 26240
rect 17880 26200 18052 26228
rect 18046 26188 18052 26200
rect 18104 26188 18110 26240
rect 21177 26231 21235 26237
rect 21177 26197 21189 26231
rect 21223 26228 21235 26231
rect 21634 26228 21640 26240
rect 21223 26200 21640 26228
rect 21223 26197 21235 26200
rect 21177 26191 21235 26197
rect 21634 26188 21640 26200
rect 21692 26188 21698 26240
rect 1104 26138 26864 26160
rect 1104 26086 3658 26138
rect 3710 26086 3722 26138
rect 3774 26086 3786 26138
rect 3838 26086 3850 26138
rect 3902 26086 3914 26138
rect 3966 26086 3978 26138
rect 4030 26086 7658 26138
rect 7710 26086 7722 26138
rect 7774 26086 7786 26138
rect 7838 26086 7850 26138
rect 7902 26086 7914 26138
rect 7966 26086 7978 26138
rect 8030 26086 11658 26138
rect 11710 26086 11722 26138
rect 11774 26086 11786 26138
rect 11838 26086 11850 26138
rect 11902 26086 11914 26138
rect 11966 26086 11978 26138
rect 12030 26086 15658 26138
rect 15710 26086 15722 26138
rect 15774 26086 15786 26138
rect 15838 26086 15850 26138
rect 15902 26086 15914 26138
rect 15966 26086 15978 26138
rect 16030 26086 19658 26138
rect 19710 26086 19722 26138
rect 19774 26086 19786 26138
rect 19838 26086 19850 26138
rect 19902 26086 19914 26138
rect 19966 26086 19978 26138
rect 20030 26086 23658 26138
rect 23710 26086 23722 26138
rect 23774 26086 23786 26138
rect 23838 26086 23850 26138
rect 23902 26086 23914 26138
rect 23966 26086 23978 26138
rect 24030 26086 26864 26138
rect 1104 26064 26864 26086
rect 4982 25984 4988 26036
rect 5040 26024 5046 26036
rect 5077 26027 5135 26033
rect 5077 26024 5089 26027
rect 5040 25996 5089 26024
rect 5040 25984 5046 25996
rect 5077 25993 5089 25996
rect 5123 25993 5135 26027
rect 5077 25987 5135 25993
rect 8389 26027 8447 26033
rect 8389 25993 8401 26027
rect 8435 26024 8447 26027
rect 9306 26024 9312 26036
rect 8435 25996 9312 26024
rect 8435 25993 8447 25996
rect 8389 25987 8447 25993
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 9585 26027 9643 26033
rect 9585 25993 9597 26027
rect 9631 26024 9643 26027
rect 9766 26024 9772 26036
rect 9631 25996 9772 26024
rect 9631 25993 9643 25996
rect 9585 25987 9643 25993
rect 9766 25984 9772 25996
rect 9824 25984 9830 26036
rect 10410 25984 10416 26036
rect 10468 26024 10474 26036
rect 15562 26024 15568 26036
rect 10468 25996 11376 26024
rect 10468 25984 10474 25996
rect 4430 25956 4436 25968
rect 3620 25928 4436 25956
rect 3620 25897 3648 25928
rect 4430 25916 4436 25928
rect 4488 25916 4494 25968
rect 5537 25959 5595 25965
rect 5537 25925 5549 25959
rect 5583 25956 5595 25959
rect 6822 25956 6828 25968
rect 5583 25928 6828 25956
rect 5583 25925 5595 25928
rect 5537 25919 5595 25925
rect 6822 25916 6828 25928
rect 6880 25916 6886 25968
rect 7098 25916 7104 25968
rect 7156 25956 7162 25968
rect 7254 25959 7312 25965
rect 7254 25956 7266 25959
rect 7156 25928 7266 25956
rect 7156 25916 7162 25928
rect 7254 25925 7266 25928
rect 7300 25925 7312 25959
rect 7254 25919 7312 25925
rect 11057 25959 11115 25965
rect 11057 25925 11069 25959
rect 11103 25956 11115 25959
rect 11146 25956 11152 25968
rect 11103 25928 11152 25956
rect 11103 25925 11115 25928
rect 11057 25919 11115 25925
rect 11146 25916 11152 25928
rect 11204 25916 11210 25968
rect 3605 25891 3663 25897
rect 3605 25857 3617 25891
rect 3651 25857 3663 25891
rect 3861 25891 3919 25897
rect 3861 25888 3873 25891
rect 3605 25851 3663 25857
rect 3712 25860 3873 25888
rect 3510 25780 3516 25832
rect 3568 25820 3574 25832
rect 3712 25820 3740 25860
rect 3861 25857 3873 25860
rect 3907 25857 3919 25891
rect 3861 25851 3919 25857
rect 5074 25848 5080 25900
rect 5132 25888 5138 25900
rect 5445 25891 5503 25897
rect 5445 25888 5457 25891
rect 5132 25860 5457 25888
rect 5132 25848 5138 25860
rect 5445 25857 5457 25860
rect 5491 25857 5503 25891
rect 5445 25851 5503 25857
rect 6086 25848 6092 25900
rect 6144 25848 6150 25900
rect 7006 25848 7012 25900
rect 7064 25848 7070 25900
rect 9030 25848 9036 25900
rect 9088 25848 9094 25900
rect 9309 25891 9367 25897
rect 9309 25857 9321 25891
rect 9355 25857 9367 25891
rect 9309 25851 9367 25857
rect 3568 25792 3740 25820
rect 3568 25780 3574 25792
rect 4982 25780 4988 25832
rect 5040 25820 5046 25832
rect 5629 25823 5687 25829
rect 5629 25820 5641 25823
rect 5040 25792 5641 25820
rect 5040 25780 5046 25792
rect 5629 25789 5641 25792
rect 5675 25789 5687 25823
rect 5629 25783 5687 25789
rect 9324 25752 9352 25851
rect 9968 25820 9996 25874
rect 11348 25829 11376 25996
rect 13004 25996 15568 26024
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25888 11759 25891
rect 12250 25888 12256 25900
rect 11747 25860 12256 25888
rect 11747 25857 11759 25860
rect 11701 25851 11759 25857
rect 12250 25848 12256 25860
rect 12308 25848 12314 25900
rect 13004 25829 13032 25996
rect 15562 25984 15568 25996
rect 15620 26024 15626 26036
rect 16666 26024 16672 26036
rect 15620 25996 16672 26024
rect 15620 25984 15626 25996
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 17129 26027 17187 26033
rect 17129 25993 17141 26027
rect 17175 26024 17187 26027
rect 17310 26024 17316 26036
rect 17175 25996 17316 26024
rect 17175 25993 17187 25996
rect 17129 25987 17187 25993
rect 17310 25984 17316 25996
rect 17368 25984 17374 26036
rect 17678 25984 17684 26036
rect 17736 26024 17742 26036
rect 17736 25996 17816 26024
rect 17736 25984 17742 25996
rect 13265 25959 13323 25965
rect 13265 25925 13277 25959
rect 13311 25956 13323 25959
rect 13354 25956 13360 25968
rect 13311 25928 13360 25956
rect 13311 25925 13323 25928
rect 13265 25919 13323 25925
rect 13354 25916 13360 25928
rect 13412 25916 13418 25968
rect 14642 25956 14648 25968
rect 14490 25928 14648 25956
rect 14642 25916 14648 25928
rect 14700 25916 14706 25968
rect 15188 25959 15246 25965
rect 15188 25925 15200 25959
rect 15234 25956 15246 25959
rect 15378 25956 15384 25968
rect 15234 25928 15384 25956
rect 15234 25925 15246 25928
rect 15188 25919 15246 25925
rect 15378 25916 15384 25928
rect 15436 25916 15442 25968
rect 17788 25965 17816 25996
rect 18046 25984 18052 26036
rect 18104 25984 18110 26036
rect 18598 25984 18604 26036
rect 18656 26024 18662 26036
rect 18785 26027 18843 26033
rect 18785 26024 18797 26027
rect 18656 25996 18797 26024
rect 18656 25984 18662 25996
rect 18785 25993 18797 25996
rect 18831 25993 18843 26027
rect 18785 25987 18843 25993
rect 18877 26027 18935 26033
rect 18877 25993 18889 26027
rect 18923 25993 18935 26027
rect 18877 25987 18935 25993
rect 19245 26027 19303 26033
rect 19245 25993 19257 26027
rect 19291 26024 19303 26027
rect 20070 26024 20076 26036
rect 19291 25996 20076 26024
rect 19291 25993 19303 25996
rect 19245 25987 19303 25993
rect 17773 25959 17831 25965
rect 17773 25925 17785 25959
rect 17819 25925 17831 25959
rect 17773 25919 17831 25925
rect 16114 25848 16120 25900
rect 16172 25888 16178 25900
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 16172 25860 17049 25888
rect 16172 25848 16178 25860
rect 17037 25857 17049 25860
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 17494 25848 17500 25900
rect 17552 25848 17558 25900
rect 17678 25848 17684 25900
rect 17736 25848 17742 25900
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25888 17923 25891
rect 18046 25888 18052 25900
rect 17911 25860 18052 25888
rect 17911 25857 17923 25860
rect 17865 25851 17923 25857
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25888 18659 25891
rect 18892 25888 18920 25987
rect 20070 25984 20076 25996
rect 20128 25984 20134 26036
rect 22646 25984 22652 26036
rect 22704 25984 22710 26036
rect 21913 25959 21971 25965
rect 21913 25956 21925 25959
rect 20930 25928 21925 25956
rect 21913 25925 21925 25928
rect 21959 25925 21971 25959
rect 22094 25956 22100 25968
rect 21913 25919 21971 25925
rect 22020 25928 22100 25956
rect 22020 25897 22048 25928
rect 22094 25916 22100 25928
rect 22152 25956 22158 25968
rect 22664 25956 22692 25984
rect 22152 25928 22692 25956
rect 22152 25916 22158 25928
rect 23474 25916 23480 25968
rect 23532 25916 23538 25968
rect 18647 25860 18920 25888
rect 22005 25891 22063 25897
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 22005 25857 22017 25891
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 11333 25823 11391 25829
rect 9968 25792 11284 25820
rect 9674 25752 9680 25764
rect 9324 25724 9680 25752
rect 9674 25712 9680 25724
rect 9732 25752 9738 25764
rect 9950 25752 9956 25764
rect 9732 25724 9956 25752
rect 9732 25712 9738 25724
rect 9950 25712 9956 25724
rect 10008 25712 10014 25764
rect 11256 25752 11284 25792
rect 11333 25789 11345 25823
rect 11379 25820 11391 25823
rect 12989 25823 13047 25829
rect 12989 25820 13001 25823
rect 11379 25792 13001 25820
rect 11379 25789 11391 25792
rect 11333 25783 11391 25789
rect 12989 25789 13001 25792
rect 13035 25789 13047 25823
rect 12989 25783 13047 25789
rect 14274 25780 14280 25832
rect 14332 25820 14338 25832
rect 14921 25823 14979 25829
rect 14921 25820 14933 25823
rect 14332 25792 14933 25820
rect 14332 25780 14338 25792
rect 14921 25789 14933 25792
rect 14967 25789 14979 25823
rect 14921 25783 14979 25789
rect 17218 25780 17224 25832
rect 17276 25780 17282 25832
rect 19337 25823 19395 25829
rect 19337 25820 19349 25823
rect 17328 25792 19349 25820
rect 11609 25755 11667 25761
rect 11609 25752 11621 25755
rect 11256 25724 11621 25752
rect 11609 25721 11621 25724
rect 11655 25721 11667 25755
rect 11609 25715 11667 25721
rect 14458 25712 14464 25764
rect 14516 25752 14522 25764
rect 14737 25755 14795 25761
rect 14737 25752 14749 25755
rect 14516 25724 14749 25752
rect 14516 25712 14522 25724
rect 14737 25721 14749 25724
rect 14783 25721 14795 25755
rect 14737 25715 14795 25721
rect 16574 25712 16580 25764
rect 16632 25752 16638 25764
rect 16669 25755 16727 25761
rect 16669 25752 16681 25755
rect 16632 25724 16681 25752
rect 16632 25712 16638 25724
rect 16669 25721 16681 25724
rect 16715 25721 16727 25755
rect 16669 25715 16727 25721
rect 4985 25687 5043 25693
rect 4985 25653 4997 25687
rect 5031 25684 5043 25687
rect 5166 25684 5172 25696
rect 5031 25656 5172 25684
rect 5031 25653 5043 25656
rect 4985 25647 5043 25653
rect 5166 25644 5172 25656
rect 5224 25644 5230 25696
rect 5902 25644 5908 25696
rect 5960 25644 5966 25696
rect 9125 25687 9183 25693
rect 9125 25653 9137 25687
rect 9171 25684 9183 25687
rect 9214 25684 9220 25696
rect 9171 25656 9220 25684
rect 9171 25653 9183 25656
rect 9125 25647 9183 25653
rect 9214 25644 9220 25656
rect 9272 25644 9278 25696
rect 9493 25687 9551 25693
rect 9493 25653 9505 25687
rect 9539 25684 9551 25687
rect 10686 25684 10692 25696
rect 9539 25656 10692 25684
rect 9539 25653 9551 25656
rect 9493 25647 9551 25653
rect 10686 25644 10692 25656
rect 10744 25644 10750 25696
rect 16298 25644 16304 25696
rect 16356 25644 16362 25696
rect 16390 25644 16396 25696
rect 16448 25684 16454 25696
rect 17328 25684 17356 25792
rect 19337 25789 19349 25792
rect 19383 25789 19395 25823
rect 19337 25783 19395 25789
rect 19429 25823 19487 25829
rect 19429 25789 19441 25823
rect 19475 25789 19487 25823
rect 19429 25783 19487 25789
rect 17862 25712 17868 25764
rect 17920 25752 17926 25764
rect 18230 25752 18236 25764
rect 17920 25724 18236 25752
rect 17920 25712 17926 25724
rect 18230 25712 18236 25724
rect 18288 25752 18294 25764
rect 19444 25752 19472 25783
rect 21358 25780 21364 25832
rect 21416 25780 21422 25832
rect 21637 25823 21695 25829
rect 21637 25789 21649 25823
rect 21683 25820 21695 25823
rect 22094 25820 22100 25832
rect 21683 25792 22100 25820
rect 21683 25789 21695 25792
rect 21637 25783 21695 25789
rect 22094 25780 22100 25792
rect 22152 25820 22158 25832
rect 22189 25823 22247 25829
rect 22189 25820 22201 25823
rect 22152 25792 22201 25820
rect 22152 25780 22158 25792
rect 22189 25789 22201 25792
rect 22235 25789 22247 25823
rect 22189 25783 22247 25789
rect 22462 25780 22468 25832
rect 22520 25780 22526 25832
rect 24213 25823 24271 25829
rect 24213 25789 24225 25823
rect 24259 25789 24271 25823
rect 24213 25783 24271 25789
rect 18288 25724 19472 25752
rect 18288 25712 18294 25724
rect 23566 25712 23572 25764
rect 23624 25752 23630 25764
rect 24228 25752 24256 25783
rect 23624 25724 24256 25752
rect 23624 25712 23630 25724
rect 16448 25656 17356 25684
rect 16448 25644 16454 25656
rect 19334 25644 19340 25696
rect 19392 25684 19398 25696
rect 19889 25687 19947 25693
rect 19889 25684 19901 25687
rect 19392 25656 19901 25684
rect 19392 25644 19398 25656
rect 19889 25653 19901 25656
rect 19935 25653 19947 25687
rect 19889 25647 19947 25653
rect 1104 25594 26864 25616
rect 1104 25542 2918 25594
rect 2970 25542 2982 25594
rect 3034 25542 3046 25594
rect 3098 25542 3110 25594
rect 3162 25542 3174 25594
rect 3226 25542 3238 25594
rect 3290 25542 6918 25594
rect 6970 25542 6982 25594
rect 7034 25542 7046 25594
rect 7098 25542 7110 25594
rect 7162 25542 7174 25594
rect 7226 25542 7238 25594
rect 7290 25542 10918 25594
rect 10970 25542 10982 25594
rect 11034 25542 11046 25594
rect 11098 25542 11110 25594
rect 11162 25542 11174 25594
rect 11226 25542 11238 25594
rect 11290 25542 14918 25594
rect 14970 25542 14982 25594
rect 15034 25542 15046 25594
rect 15098 25542 15110 25594
rect 15162 25542 15174 25594
rect 15226 25542 15238 25594
rect 15290 25542 18918 25594
rect 18970 25542 18982 25594
rect 19034 25542 19046 25594
rect 19098 25542 19110 25594
rect 19162 25542 19174 25594
rect 19226 25542 19238 25594
rect 19290 25542 22918 25594
rect 22970 25542 22982 25594
rect 23034 25542 23046 25594
rect 23098 25542 23110 25594
rect 23162 25542 23174 25594
rect 23226 25542 23238 25594
rect 23290 25542 26864 25594
rect 1104 25520 26864 25542
rect 4062 25440 4068 25492
rect 4120 25440 4126 25492
rect 12986 25440 12992 25492
rect 13044 25440 13050 25492
rect 15289 25483 15347 25489
rect 15289 25449 15301 25483
rect 15335 25480 15347 25483
rect 15378 25480 15384 25492
rect 15335 25452 15384 25480
rect 15335 25449 15347 25452
rect 15289 25443 15347 25449
rect 15378 25440 15384 25452
rect 15436 25440 15442 25492
rect 17405 25483 17463 25489
rect 17405 25449 17417 25483
rect 17451 25480 17463 25483
rect 17954 25480 17960 25492
rect 17451 25452 17960 25480
rect 17451 25449 17463 25452
rect 17405 25443 17463 25449
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 19518 25440 19524 25492
rect 19576 25480 19582 25492
rect 19797 25483 19855 25489
rect 19797 25480 19809 25483
rect 19576 25452 19809 25480
rect 19576 25440 19582 25452
rect 19797 25449 19809 25452
rect 19843 25449 19855 25483
rect 19797 25443 19855 25449
rect 8757 25415 8815 25421
rect 8757 25381 8769 25415
rect 8803 25381 8815 25415
rect 17862 25412 17868 25424
rect 8757 25375 8815 25381
rect 13648 25384 17868 25412
rect 4709 25347 4767 25353
rect 4709 25313 4721 25347
rect 4755 25344 4767 25347
rect 4982 25344 4988 25356
rect 4755 25316 4988 25344
rect 4755 25313 4767 25316
rect 4709 25307 4767 25313
rect 4982 25304 4988 25316
rect 5040 25304 5046 25356
rect 7374 25304 7380 25356
rect 7432 25304 7438 25356
rect 8772 25344 8800 25375
rect 8846 25344 8852 25356
rect 8772 25316 8852 25344
rect 8846 25304 8852 25316
rect 8904 25344 8910 25356
rect 9585 25347 9643 25353
rect 9585 25344 9597 25347
rect 8904 25316 9597 25344
rect 8904 25304 8910 25316
rect 9585 25313 9597 25316
rect 9631 25313 9643 25347
rect 9585 25307 9643 25313
rect 12342 25304 12348 25356
rect 12400 25344 12406 25356
rect 13648 25353 13676 25384
rect 17862 25372 17868 25384
rect 17920 25372 17926 25424
rect 22097 25415 22155 25421
rect 22097 25381 22109 25415
rect 22143 25412 22155 25415
rect 22462 25412 22468 25424
rect 22143 25384 22468 25412
rect 22143 25381 22155 25384
rect 22097 25375 22155 25381
rect 22462 25372 22468 25384
rect 22520 25372 22526 25424
rect 13633 25347 13691 25353
rect 13633 25344 13645 25347
rect 12400 25316 13645 25344
rect 12400 25304 12406 25316
rect 13633 25313 13645 25316
rect 13679 25313 13691 25347
rect 13633 25307 13691 25313
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25344 16175 25347
rect 16482 25344 16488 25356
rect 16163 25316 16488 25344
rect 16163 25313 16175 25316
rect 16117 25307 16175 25313
rect 16482 25304 16488 25316
rect 16540 25304 16546 25356
rect 18046 25304 18052 25356
rect 18104 25344 18110 25356
rect 21174 25344 21180 25356
rect 18104 25316 21180 25344
rect 18104 25304 18110 25316
rect 5353 25279 5411 25285
rect 5353 25245 5365 25279
rect 5399 25276 5411 25279
rect 5442 25276 5448 25288
rect 5399 25248 5448 25276
rect 5399 25245 5411 25248
rect 5353 25239 5411 25245
rect 5442 25236 5448 25248
rect 5500 25236 5506 25288
rect 5620 25279 5678 25285
rect 5620 25245 5632 25279
rect 5666 25276 5678 25279
rect 5902 25276 5908 25288
rect 5666 25248 5908 25276
rect 5666 25245 5678 25248
rect 5620 25239 5678 25245
rect 5902 25236 5908 25248
rect 5960 25236 5966 25288
rect 9122 25236 9128 25288
rect 9180 25236 9186 25288
rect 9214 25236 9220 25288
rect 9272 25276 9278 25288
rect 9677 25279 9735 25285
rect 9677 25276 9689 25279
rect 9272 25248 9689 25276
rect 9272 25236 9278 25248
rect 9677 25245 9689 25248
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 9861 25279 9919 25285
rect 9861 25245 9873 25279
rect 9907 25276 9919 25279
rect 9950 25276 9956 25288
rect 9907 25248 9956 25276
rect 9907 25245 9919 25248
rect 9861 25239 9919 25245
rect 9950 25236 9956 25248
rect 10008 25236 10014 25288
rect 10229 25279 10287 25285
rect 10229 25245 10241 25279
rect 10275 25245 10287 25279
rect 10229 25239 10287 25245
rect 4433 25211 4491 25217
rect 4433 25177 4445 25211
rect 4479 25208 4491 25211
rect 5166 25208 5172 25220
rect 4479 25180 5172 25208
rect 4479 25177 4491 25180
rect 4433 25171 4491 25177
rect 5166 25168 5172 25180
rect 5224 25168 5230 25220
rect 7644 25211 7702 25217
rect 7644 25177 7656 25211
rect 7690 25208 7702 25211
rect 10244 25208 10272 25239
rect 12250 25236 12256 25288
rect 12308 25236 12314 25288
rect 13357 25279 13415 25285
rect 13357 25245 13369 25279
rect 13403 25276 13415 25279
rect 13814 25276 13820 25288
rect 13403 25248 13820 25276
rect 13403 25245 13415 25248
rect 13357 25239 13415 25245
rect 13814 25236 13820 25248
rect 13872 25236 13878 25288
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25276 15531 25279
rect 17221 25279 17279 25285
rect 15519 25248 15608 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 10410 25208 10416 25220
rect 7690 25180 8984 25208
rect 10244 25180 10416 25208
rect 7690 25177 7702 25180
rect 7644 25171 7702 25177
rect 4525 25143 4583 25149
rect 4525 25109 4537 25143
rect 4571 25140 4583 25143
rect 5902 25140 5908 25152
rect 4571 25112 5908 25140
rect 4571 25109 4583 25112
rect 4525 25103 4583 25109
rect 5902 25100 5908 25112
rect 5960 25140 5966 25152
rect 6454 25140 6460 25152
rect 5960 25112 6460 25140
rect 5960 25100 5966 25112
rect 6454 25100 6460 25112
rect 6512 25100 6518 25152
rect 6546 25100 6552 25152
rect 6604 25140 6610 25152
rect 8956 25149 8984 25180
rect 10410 25168 10416 25180
rect 10468 25168 10474 25220
rect 10502 25168 10508 25220
rect 10560 25168 10566 25220
rect 12161 25211 12219 25217
rect 12161 25208 12173 25211
rect 11730 25180 12173 25208
rect 12161 25177 12173 25180
rect 12207 25177 12219 25211
rect 12161 25171 12219 25177
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 6604 25112 6745 25140
rect 6604 25100 6610 25112
rect 6733 25109 6745 25112
rect 6779 25109 6791 25143
rect 6733 25103 6791 25109
rect 8941 25143 8999 25149
rect 8941 25109 8953 25143
rect 8987 25109 8999 25143
rect 8941 25103 8999 25109
rect 10045 25143 10103 25149
rect 10045 25109 10057 25143
rect 10091 25140 10103 25143
rect 10318 25140 10324 25152
rect 10091 25112 10324 25140
rect 10091 25109 10103 25112
rect 10045 25103 10103 25109
rect 10318 25100 10324 25112
rect 10376 25100 10382 25152
rect 11514 25100 11520 25152
rect 11572 25140 11578 25152
rect 11977 25143 12035 25149
rect 11977 25140 11989 25143
rect 11572 25112 11989 25140
rect 11572 25100 11578 25112
rect 11977 25109 11989 25112
rect 12023 25109 12035 25143
rect 11977 25103 12035 25109
rect 13446 25100 13452 25152
rect 13504 25100 13510 25152
rect 15580 25149 15608 25248
rect 17221 25245 17233 25279
rect 17267 25276 17279 25279
rect 17402 25276 17408 25288
rect 17267 25248 17408 25276
rect 17267 25245 17279 25248
rect 17221 25239 17279 25245
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 19628 25285 19656 25316
rect 21174 25304 21180 25316
rect 21232 25304 21238 25356
rect 21634 25304 21640 25356
rect 21692 25304 21698 25356
rect 23566 25344 23572 25356
rect 21744 25316 23572 25344
rect 21744 25285 21772 25316
rect 23566 25304 23572 25316
rect 23624 25304 23630 25356
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 18748 25248 19257 25276
rect 18748 25236 18754 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 21085 25279 21143 25285
rect 21085 25245 21097 25279
rect 21131 25245 21143 25279
rect 21085 25239 21143 25245
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25245 21787 25279
rect 21729 25239 21787 25245
rect 15933 25211 15991 25217
rect 15933 25177 15945 25211
rect 15979 25208 15991 25211
rect 16298 25208 16304 25220
rect 15979 25180 16304 25208
rect 15979 25177 15991 25180
rect 15933 25171 15991 25177
rect 16298 25168 16304 25180
rect 16356 25168 16362 25220
rect 19429 25211 19487 25217
rect 19429 25177 19441 25211
rect 19475 25177 19487 25211
rect 19429 25171 19487 25177
rect 19521 25211 19579 25217
rect 19521 25177 19533 25211
rect 19567 25208 19579 25211
rect 20530 25208 20536 25220
rect 19567 25180 20536 25208
rect 19567 25177 19579 25180
rect 19521 25171 19579 25177
rect 15565 25143 15623 25149
rect 15565 25109 15577 25143
rect 15611 25109 15623 25143
rect 15565 25103 15623 25109
rect 16025 25143 16083 25149
rect 16025 25109 16037 25143
rect 16071 25140 16083 25143
rect 16206 25140 16212 25152
rect 16071 25112 16212 25140
rect 16071 25109 16083 25112
rect 16025 25103 16083 25109
rect 16206 25100 16212 25112
rect 16264 25140 16270 25152
rect 17310 25140 17316 25152
rect 16264 25112 17316 25140
rect 16264 25100 16270 25112
rect 17310 25100 17316 25112
rect 17368 25100 17374 25152
rect 19444 25140 19472 25171
rect 20530 25168 20536 25180
rect 20588 25168 20594 25220
rect 20806 25168 20812 25220
rect 20864 25168 20870 25220
rect 21100 25208 21128 25239
rect 22554 25236 22560 25288
rect 22612 25276 22618 25288
rect 22925 25279 22983 25285
rect 22925 25276 22937 25279
rect 22612 25248 22937 25276
rect 22612 25236 22618 25248
rect 22925 25245 22937 25248
rect 22971 25245 22983 25279
rect 22925 25239 22983 25245
rect 21100 25180 22692 25208
rect 22664 25152 22692 25180
rect 20622 25140 20628 25152
rect 19444 25112 20628 25140
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 22646 25100 22652 25152
rect 22704 25140 22710 25152
rect 23017 25143 23075 25149
rect 23017 25140 23029 25143
rect 22704 25112 23029 25140
rect 22704 25100 22710 25112
rect 23017 25109 23029 25112
rect 23063 25109 23075 25143
rect 23017 25103 23075 25109
rect 1104 25050 26864 25072
rect 1104 24998 3658 25050
rect 3710 24998 3722 25050
rect 3774 24998 3786 25050
rect 3838 24998 3850 25050
rect 3902 24998 3914 25050
rect 3966 24998 3978 25050
rect 4030 24998 7658 25050
rect 7710 24998 7722 25050
rect 7774 24998 7786 25050
rect 7838 24998 7850 25050
rect 7902 24998 7914 25050
rect 7966 24998 7978 25050
rect 8030 24998 11658 25050
rect 11710 24998 11722 25050
rect 11774 24998 11786 25050
rect 11838 24998 11850 25050
rect 11902 24998 11914 25050
rect 11966 24998 11978 25050
rect 12030 24998 15658 25050
rect 15710 24998 15722 25050
rect 15774 24998 15786 25050
rect 15838 24998 15850 25050
rect 15902 24998 15914 25050
rect 15966 24998 15978 25050
rect 16030 24998 19658 25050
rect 19710 24998 19722 25050
rect 19774 24998 19786 25050
rect 19838 24998 19850 25050
rect 19902 24998 19914 25050
rect 19966 24998 19978 25050
rect 20030 24998 23658 25050
rect 23710 24998 23722 25050
rect 23774 24998 23786 25050
rect 23838 24998 23850 25050
rect 23902 24998 23914 25050
rect 23966 24998 23978 25050
rect 24030 24998 26864 25050
rect 1104 24976 26864 24998
rect 6086 24896 6092 24948
rect 6144 24936 6150 24948
rect 6365 24939 6423 24945
rect 6365 24936 6377 24939
rect 6144 24908 6377 24936
rect 6144 24896 6150 24908
rect 6365 24905 6377 24908
rect 6411 24905 6423 24939
rect 6365 24899 6423 24905
rect 6454 24896 6460 24948
rect 6512 24936 6518 24948
rect 6512 24908 6868 24936
rect 6512 24896 6518 24908
rect 6546 24828 6552 24880
rect 6604 24868 6610 24880
rect 6840 24877 6868 24908
rect 8846 24896 8852 24948
rect 8904 24896 8910 24948
rect 9122 24896 9128 24948
rect 9180 24936 9186 24948
rect 9217 24939 9275 24945
rect 9217 24936 9229 24939
rect 9180 24908 9229 24936
rect 9180 24896 9186 24908
rect 9217 24905 9229 24908
rect 9263 24905 9275 24939
rect 9217 24899 9275 24905
rect 10502 24896 10508 24948
rect 10560 24936 10566 24948
rect 10873 24939 10931 24945
rect 10873 24936 10885 24939
rect 10560 24908 10885 24936
rect 10560 24896 10566 24908
rect 10873 24905 10885 24908
rect 10919 24905 10931 24939
rect 10873 24899 10931 24905
rect 15562 24896 15568 24948
rect 15620 24936 15626 24948
rect 18046 24936 18052 24948
rect 15620 24908 18052 24936
rect 15620 24896 15626 24908
rect 18046 24896 18052 24908
rect 18104 24896 18110 24948
rect 6733 24871 6791 24877
rect 6733 24868 6745 24871
rect 6604 24840 6745 24868
rect 6604 24828 6610 24840
rect 6733 24837 6745 24840
rect 6779 24837 6791 24871
rect 6733 24831 6791 24837
rect 6825 24871 6883 24877
rect 6825 24837 6837 24871
rect 6871 24868 6883 24871
rect 9398 24868 9404 24880
rect 6871 24840 9404 24868
rect 6871 24837 6883 24840
rect 6825 24831 6883 24837
rect 9398 24828 9404 24840
rect 9456 24828 9462 24880
rect 2501 24803 2559 24809
rect 2501 24769 2513 24803
rect 2547 24800 2559 24803
rect 3053 24803 3111 24809
rect 2547 24772 2728 24800
rect 2547 24769 2559 24772
rect 2501 24763 2559 24769
rect 2700 24673 2728 24772
rect 3053 24769 3065 24803
rect 3099 24800 3111 24803
rect 3510 24800 3516 24812
rect 3099 24772 3516 24800
rect 3099 24769 3111 24772
rect 3053 24763 3111 24769
rect 3510 24760 3516 24772
rect 3568 24760 3574 24812
rect 5350 24760 5356 24812
rect 5408 24800 5414 24812
rect 5445 24803 5503 24809
rect 5445 24800 5457 24803
rect 5408 24772 5457 24800
rect 5408 24760 5414 24772
rect 5445 24769 5457 24772
rect 5491 24769 5503 24803
rect 8757 24803 8815 24809
rect 8757 24800 8769 24803
rect 5445 24763 5503 24769
rect 5552 24772 8769 24800
rect 3145 24735 3203 24741
rect 3145 24701 3157 24735
rect 3191 24701 3203 24735
rect 3145 24695 3203 24701
rect 3329 24735 3387 24741
rect 3329 24701 3341 24735
rect 3375 24732 3387 24735
rect 4982 24732 4988 24744
rect 3375 24704 4988 24732
rect 3375 24701 3387 24704
rect 3329 24695 3387 24701
rect 2685 24667 2743 24673
rect 2685 24633 2697 24667
rect 2731 24633 2743 24667
rect 3160 24664 3188 24695
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 4062 24664 4068 24676
rect 3160 24636 4068 24664
rect 2685 24627 2743 24633
rect 3344 24608 3372 24636
rect 4062 24624 4068 24636
rect 4120 24664 4126 24676
rect 5552 24664 5580 24772
rect 8757 24769 8769 24772
rect 8803 24769 8815 24803
rect 8757 24763 8815 24769
rect 10318 24760 10324 24812
rect 10376 24760 10382 24812
rect 10502 24760 10508 24812
rect 10560 24760 10566 24812
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24732 7067 24735
rect 7558 24732 7564 24744
rect 7055 24704 7564 24732
rect 7055 24701 7067 24704
rect 7009 24695 7067 24701
rect 7558 24692 7564 24704
rect 7616 24692 7622 24744
rect 8662 24692 8668 24744
rect 8720 24732 8726 24744
rect 8938 24732 8944 24744
rect 8720 24704 8944 24732
rect 8720 24692 8726 24704
rect 8938 24692 8944 24704
rect 8996 24692 9002 24744
rect 10612 24732 10640 24763
rect 10686 24760 10692 24812
rect 10744 24760 10750 24812
rect 13538 24760 13544 24812
rect 13596 24800 13602 24812
rect 15562 24800 15568 24812
rect 13596 24772 15568 24800
rect 13596 24760 13602 24772
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 19153 24803 19211 24809
rect 19153 24769 19165 24803
rect 19199 24800 19211 24803
rect 19334 24800 19340 24812
rect 19199 24772 19340 24800
rect 19199 24769 19211 24772
rect 19153 24763 19211 24769
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 19518 24760 19524 24812
rect 19576 24800 19582 24812
rect 19797 24803 19855 24809
rect 19797 24800 19809 24803
rect 19576 24772 19809 24800
rect 19576 24760 19582 24772
rect 19797 24769 19809 24772
rect 19843 24769 19855 24803
rect 19797 24763 19855 24769
rect 11514 24732 11520 24744
rect 10612 24704 11520 24732
rect 11514 24692 11520 24704
rect 11572 24692 11578 24744
rect 19886 24692 19892 24744
rect 19944 24692 19950 24744
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24732 20223 24735
rect 21358 24732 21364 24744
rect 20211 24704 21364 24732
rect 20211 24701 20223 24704
rect 20165 24695 20223 24701
rect 21358 24692 21364 24704
rect 21416 24692 21422 24744
rect 4120 24636 5580 24664
rect 4120 24624 4126 24636
rect 10318 24624 10324 24676
rect 10376 24664 10382 24676
rect 10686 24664 10692 24676
rect 10376 24636 10692 24664
rect 10376 24624 10382 24636
rect 10686 24624 10692 24636
rect 10744 24624 10750 24676
rect 2130 24556 2136 24608
rect 2188 24596 2194 24608
rect 2317 24599 2375 24605
rect 2317 24596 2329 24599
rect 2188 24568 2329 24596
rect 2188 24556 2194 24568
rect 2317 24565 2329 24568
rect 2363 24565 2375 24599
rect 2317 24559 2375 24565
rect 3326 24556 3332 24608
rect 3384 24556 3390 24608
rect 5258 24556 5264 24608
rect 5316 24556 5322 24608
rect 19429 24599 19487 24605
rect 19429 24565 19441 24599
rect 19475 24596 19487 24599
rect 19518 24596 19524 24608
rect 19475 24568 19524 24596
rect 19475 24565 19487 24568
rect 19429 24559 19487 24565
rect 19518 24556 19524 24568
rect 19576 24556 19582 24608
rect 1104 24506 26864 24528
rect 1104 24454 2918 24506
rect 2970 24454 2982 24506
rect 3034 24454 3046 24506
rect 3098 24454 3110 24506
rect 3162 24454 3174 24506
rect 3226 24454 3238 24506
rect 3290 24454 6918 24506
rect 6970 24454 6982 24506
rect 7034 24454 7046 24506
rect 7098 24454 7110 24506
rect 7162 24454 7174 24506
rect 7226 24454 7238 24506
rect 7290 24454 10918 24506
rect 10970 24454 10982 24506
rect 11034 24454 11046 24506
rect 11098 24454 11110 24506
rect 11162 24454 11174 24506
rect 11226 24454 11238 24506
rect 11290 24454 14918 24506
rect 14970 24454 14982 24506
rect 15034 24454 15046 24506
rect 15098 24454 15110 24506
rect 15162 24454 15174 24506
rect 15226 24454 15238 24506
rect 15290 24454 18918 24506
rect 18970 24454 18982 24506
rect 19034 24454 19046 24506
rect 19098 24454 19110 24506
rect 19162 24454 19174 24506
rect 19226 24454 19238 24506
rect 19290 24454 22918 24506
rect 22970 24454 22982 24506
rect 23034 24454 23046 24506
rect 23098 24454 23110 24506
rect 23162 24454 23174 24506
rect 23226 24454 23238 24506
rect 23290 24454 26864 24506
rect 1104 24432 26864 24454
rect 23474 24216 23480 24268
rect 23532 24256 23538 24268
rect 23845 24259 23903 24265
rect 23845 24256 23857 24259
rect 23532 24228 23857 24256
rect 23532 24216 23538 24228
rect 23845 24225 23857 24228
rect 23891 24225 23903 24259
rect 23845 24219 23903 24225
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 1946 24188 1952 24200
rect 1903 24160 1952 24188
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 1946 24148 1952 24160
rect 2004 24148 2010 24200
rect 2130 24197 2136 24200
rect 2124 24188 2136 24197
rect 2091 24160 2136 24188
rect 2124 24151 2136 24160
rect 2130 24148 2136 24151
rect 2188 24148 2194 24200
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24188 4951 24191
rect 5442 24188 5448 24200
rect 4939 24160 5448 24188
rect 4939 24157 4951 24160
rect 4893 24151 4951 24157
rect 4338 24080 4344 24132
rect 4396 24120 4402 24132
rect 4908 24120 4936 24151
rect 5442 24148 5448 24160
rect 5500 24148 5506 24200
rect 13354 24148 13360 24200
rect 13412 24148 13418 24200
rect 19886 24148 19892 24200
rect 19944 24148 19950 24200
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 20162 24148 20168 24200
rect 20220 24148 20226 24200
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22646 24188 22652 24200
rect 22235 24160 22652 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 22646 24148 22652 24160
rect 22704 24188 22710 24200
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 22704 24160 24409 24188
rect 22704 24148 22710 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24397 24151 24455 24157
rect 4396 24092 4936 24120
rect 5160 24123 5218 24129
rect 4396 24080 4402 24092
rect 5160 24089 5172 24123
rect 5206 24120 5218 24123
rect 5258 24120 5264 24132
rect 5206 24092 5264 24120
rect 5206 24089 5218 24092
rect 5160 24083 5218 24089
rect 5258 24080 5264 24092
rect 5316 24080 5322 24132
rect 7558 24080 7564 24132
rect 7616 24120 7622 24132
rect 13538 24120 13544 24132
rect 7616 24092 13544 24120
rect 7616 24080 7622 24092
rect 13538 24080 13544 24092
rect 13596 24080 13602 24132
rect 3237 24055 3295 24061
rect 3237 24021 3249 24055
rect 3283 24052 3295 24055
rect 3510 24052 3516 24064
rect 3283 24024 3516 24052
rect 3283 24021 3295 24024
rect 3237 24015 3295 24021
rect 3510 24012 3516 24024
rect 3568 24012 3574 24064
rect 4614 24012 4620 24064
rect 4672 24012 4678 24064
rect 6270 24012 6276 24064
rect 6328 24012 6334 24064
rect 13170 24012 13176 24064
rect 13228 24012 13234 24064
rect 19904 24052 19932 24148
rect 19981 24123 20039 24129
rect 19981 24089 19993 24123
rect 20027 24120 20039 24123
rect 20441 24123 20499 24129
rect 20441 24120 20453 24123
rect 20027 24092 20453 24120
rect 20027 24089 20039 24092
rect 19981 24083 20039 24089
rect 20441 24089 20453 24092
rect 20487 24089 20499 24123
rect 22097 24123 22155 24129
rect 22097 24120 22109 24123
rect 21666 24092 22109 24120
rect 20441 24083 20499 24089
rect 22097 24089 22109 24092
rect 22143 24089 22155 24123
rect 22097 24083 22155 24089
rect 22830 24080 22836 24132
rect 22888 24120 22894 24132
rect 23753 24123 23811 24129
rect 23753 24120 23765 24123
rect 22888 24092 23765 24120
rect 22888 24080 22894 24092
rect 23753 24089 23765 24092
rect 23799 24089 23811 24123
rect 25130 24120 25136 24132
rect 23753 24083 23811 24089
rect 24412 24092 25136 24120
rect 20254 24052 20260 24064
rect 19904 24024 20260 24052
rect 20254 24012 20260 24024
rect 20312 24012 20318 24064
rect 21358 24012 21364 24064
rect 21416 24052 21422 24064
rect 21913 24055 21971 24061
rect 21913 24052 21925 24055
rect 21416 24024 21925 24052
rect 21416 24012 21422 24024
rect 21913 24021 21925 24024
rect 21959 24021 21971 24055
rect 21913 24015 21971 24021
rect 23198 24012 23204 24064
rect 23256 24052 23262 24064
rect 23293 24055 23351 24061
rect 23293 24052 23305 24055
rect 23256 24024 23305 24052
rect 23256 24012 23262 24024
rect 23293 24021 23305 24024
rect 23339 24021 23351 24055
rect 23293 24015 23351 24021
rect 23661 24055 23719 24061
rect 23661 24021 23673 24055
rect 23707 24052 23719 24055
rect 24412 24052 24440 24092
rect 25130 24080 25136 24092
rect 25188 24080 25194 24132
rect 23707 24024 24440 24052
rect 23707 24021 23719 24024
rect 23661 24015 23719 24021
rect 24486 24012 24492 24064
rect 24544 24012 24550 24064
rect 1104 23962 26864 23984
rect 1104 23910 3658 23962
rect 3710 23910 3722 23962
rect 3774 23910 3786 23962
rect 3838 23910 3850 23962
rect 3902 23910 3914 23962
rect 3966 23910 3978 23962
rect 4030 23910 7658 23962
rect 7710 23910 7722 23962
rect 7774 23910 7786 23962
rect 7838 23910 7850 23962
rect 7902 23910 7914 23962
rect 7966 23910 7978 23962
rect 8030 23910 11658 23962
rect 11710 23910 11722 23962
rect 11774 23910 11786 23962
rect 11838 23910 11850 23962
rect 11902 23910 11914 23962
rect 11966 23910 11978 23962
rect 12030 23910 15658 23962
rect 15710 23910 15722 23962
rect 15774 23910 15786 23962
rect 15838 23910 15850 23962
rect 15902 23910 15914 23962
rect 15966 23910 15978 23962
rect 16030 23910 19658 23962
rect 19710 23910 19722 23962
rect 19774 23910 19786 23962
rect 19838 23910 19850 23962
rect 19902 23910 19914 23962
rect 19966 23910 19978 23962
rect 20030 23910 23658 23962
rect 23710 23910 23722 23962
rect 23774 23910 23786 23962
rect 23838 23910 23850 23962
rect 23902 23910 23914 23962
rect 23966 23910 23978 23962
rect 24030 23910 26864 23962
rect 1104 23888 26864 23910
rect 3513 23851 3571 23857
rect 3513 23848 3525 23851
rect 1780 23820 3525 23848
rect 1780 23721 1808 23820
rect 3513 23817 3525 23820
rect 3559 23817 3571 23851
rect 3513 23811 3571 23817
rect 3973 23851 4031 23857
rect 3973 23817 3985 23851
rect 4019 23848 4031 23851
rect 4062 23848 4068 23860
rect 4019 23820 4068 23848
rect 4019 23817 4031 23820
rect 3973 23811 4031 23817
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 4798 23808 4804 23860
rect 4856 23848 4862 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 4856 23820 6377 23848
rect 4856 23808 4862 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 6365 23811 6423 23817
rect 6822 23808 6828 23860
rect 6880 23808 6886 23860
rect 12406 23820 13308 23848
rect 4614 23789 4620 23792
rect 4608 23780 4620 23789
rect 2056 23752 4384 23780
rect 4575 23752 4620 23780
rect 1765 23715 1823 23721
rect 1765 23681 1777 23715
rect 1811 23681 1823 23715
rect 1765 23675 1823 23681
rect 1946 23672 1952 23724
rect 2004 23712 2010 23724
rect 2056 23721 2084 23752
rect 4356 23724 4384 23752
rect 4608 23743 4620 23752
rect 4614 23740 4620 23743
rect 4672 23740 4678 23792
rect 4982 23740 4988 23792
rect 5040 23780 5046 23792
rect 12406 23780 12434 23820
rect 5040 23752 12434 23780
rect 5040 23740 5046 23752
rect 12802 23740 12808 23792
rect 12860 23780 12866 23792
rect 13142 23783 13200 23789
rect 13142 23780 13154 23783
rect 12860 23752 13154 23780
rect 12860 23740 12866 23752
rect 13142 23749 13154 23752
rect 13188 23749 13200 23783
rect 13280 23780 13308 23820
rect 13446 23808 13452 23860
rect 13504 23848 13510 23860
rect 14829 23851 14887 23857
rect 14829 23848 14841 23851
rect 13504 23820 14841 23848
rect 13504 23808 13510 23820
rect 14829 23817 14841 23820
rect 14875 23817 14887 23851
rect 14829 23811 14887 23817
rect 20070 23808 20076 23860
rect 20128 23848 20134 23860
rect 20257 23851 20315 23857
rect 20257 23848 20269 23851
rect 20128 23820 20269 23848
rect 20128 23808 20134 23820
rect 20257 23817 20269 23820
rect 20303 23817 20315 23851
rect 20257 23811 20315 23817
rect 23385 23851 23443 23857
rect 23385 23817 23397 23851
rect 23431 23817 23443 23851
rect 23385 23811 23443 23817
rect 16942 23780 16948 23792
rect 13280 23752 16948 23780
rect 13142 23743 13200 23749
rect 2041 23715 2099 23721
rect 2041 23712 2053 23715
rect 2004 23684 2053 23712
rect 2004 23672 2010 23684
rect 2041 23681 2053 23684
rect 2087 23681 2099 23715
rect 2297 23715 2355 23721
rect 2297 23712 2309 23715
rect 2041 23675 2099 23681
rect 2148 23684 2309 23712
rect 2148 23644 2176 23684
rect 2297 23681 2309 23684
rect 2343 23681 2355 23715
rect 2297 23675 2355 23681
rect 3881 23715 3939 23721
rect 3881 23681 3893 23715
rect 3927 23712 3939 23715
rect 4062 23712 4068 23724
rect 3927 23684 4068 23712
rect 3927 23681 3939 23684
rect 3881 23675 3939 23681
rect 1964 23616 2176 23644
rect 1964 23585 1992 23616
rect 1949 23579 2007 23585
rect 1949 23545 1961 23579
rect 1995 23545 2007 23579
rect 1949 23539 2007 23545
rect 3421 23579 3479 23585
rect 3421 23545 3433 23579
rect 3467 23576 3479 23579
rect 3896 23576 3924 23675
rect 4062 23672 4068 23684
rect 4120 23672 4126 23724
rect 4338 23672 4344 23724
rect 4396 23672 4402 23724
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23681 6791 23715
rect 6733 23675 6791 23681
rect 4157 23647 4215 23653
rect 4157 23613 4169 23647
rect 4203 23613 4215 23647
rect 4157 23607 4215 23613
rect 3467 23548 3924 23576
rect 3467 23545 3479 23548
rect 3421 23539 3479 23545
rect 4172 23508 4200 23607
rect 5718 23536 5724 23588
rect 5776 23576 5782 23588
rect 6748 23576 6776 23675
rect 7374 23672 7380 23724
rect 7432 23712 7438 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7432 23684 7941 23712
rect 7432 23672 7438 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 11333 23715 11391 23721
rect 11333 23681 11345 23715
rect 11379 23712 11391 23715
rect 12250 23712 12256 23724
rect 11379 23684 12256 23712
rect 11379 23681 11391 23684
rect 11333 23675 11391 23681
rect 12250 23672 12256 23684
rect 12308 23672 12314 23724
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23712 12679 23715
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 12667 23684 14412 23712
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 7009 23647 7067 23653
rect 7009 23613 7021 23647
rect 7055 23644 7067 23647
rect 7466 23644 7472 23656
rect 7055 23616 7472 23644
rect 7055 23613 7067 23616
rect 7009 23607 7067 23613
rect 7466 23604 7472 23616
rect 7524 23604 7530 23656
rect 7558 23604 7564 23656
rect 7616 23644 7622 23656
rect 7653 23647 7711 23653
rect 7653 23644 7665 23647
rect 7616 23616 7665 23644
rect 7616 23604 7622 23616
rect 7653 23613 7665 23616
rect 7699 23613 7711 23647
rect 7653 23607 7711 23613
rect 7837 23647 7895 23653
rect 7837 23613 7849 23647
rect 7883 23644 7895 23647
rect 8110 23644 8116 23656
rect 7883 23616 8116 23644
rect 7883 23613 7895 23616
rect 7837 23607 7895 23613
rect 5776 23548 6776 23576
rect 5776 23536 5782 23548
rect 6822 23536 6828 23588
rect 6880 23576 6886 23588
rect 7852 23576 7880 23607
rect 8110 23604 8116 23616
rect 8168 23644 8174 23656
rect 8386 23644 8392 23656
rect 8168 23616 8392 23644
rect 8168 23604 8174 23616
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12492 23616 12909 23644
rect 12492 23604 12498 23616
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 12897 23607 12955 23613
rect 6880 23548 7880 23576
rect 6880 23536 6886 23548
rect 12802 23536 12808 23588
rect 12860 23536 12866 23588
rect 14384 23585 14412 23684
rect 14476 23684 14749 23712
rect 14369 23579 14427 23585
rect 14369 23545 14381 23579
rect 14415 23545 14427 23579
rect 14369 23539 14427 23545
rect 5994 23508 6000 23520
rect 4172 23480 6000 23508
rect 5994 23468 6000 23480
rect 6052 23468 6058 23520
rect 8297 23511 8355 23517
rect 8297 23477 8309 23511
rect 8343 23508 8355 23511
rect 8754 23508 8760 23520
rect 8343 23480 8760 23508
rect 8343 23477 8355 23480
rect 8297 23471 8355 23477
rect 8754 23468 8760 23480
rect 8812 23468 8818 23520
rect 11241 23511 11299 23517
rect 11241 23477 11253 23511
rect 11287 23508 11299 23511
rect 11330 23508 11336 23520
rect 11287 23480 11336 23508
rect 11287 23477 11299 23480
rect 11241 23471 11299 23477
rect 11330 23468 11336 23480
rect 11388 23468 11394 23520
rect 14274 23468 14280 23520
rect 14332 23508 14338 23520
rect 14476 23508 14504 23684
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 15028 23653 15056 23752
rect 16942 23740 16948 23752
rect 17000 23780 17006 23792
rect 17218 23780 17224 23792
rect 17000 23752 17224 23780
rect 17000 23740 17006 23752
rect 17218 23740 17224 23752
rect 17276 23740 17282 23792
rect 17954 23740 17960 23792
rect 18012 23740 18018 23792
rect 19153 23783 19211 23789
rect 19153 23749 19165 23783
rect 19199 23780 19211 23783
rect 19242 23780 19248 23792
rect 19199 23752 19248 23780
rect 19199 23749 19211 23752
rect 19153 23743 19211 23749
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 19337 23783 19395 23789
rect 19337 23749 19349 23783
rect 19383 23780 19395 23783
rect 19702 23780 19708 23792
rect 19383 23752 19708 23780
rect 19383 23749 19395 23752
rect 19337 23743 19395 23749
rect 19702 23740 19708 23752
rect 19760 23740 19766 23792
rect 19812 23752 20392 23780
rect 16117 23715 16175 23721
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 15013 23647 15071 23653
rect 15013 23613 15025 23647
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 15562 23604 15568 23656
rect 15620 23644 15626 23656
rect 16025 23647 16083 23653
rect 16025 23644 16037 23647
rect 15620 23616 16037 23644
rect 15620 23604 15626 23616
rect 16025 23613 16037 23616
rect 16071 23613 16083 23647
rect 16025 23607 16083 23613
rect 14332 23480 14504 23508
rect 16132 23508 16160 23675
rect 16666 23672 16672 23724
rect 16724 23672 16730 23724
rect 18414 23672 18420 23724
rect 18472 23712 18478 23724
rect 19812 23721 19840 23752
rect 19521 23715 19579 23721
rect 19521 23712 19533 23715
rect 18472 23684 19533 23712
rect 18472 23672 18478 23684
rect 19521 23681 19533 23684
rect 19567 23681 19579 23715
rect 19521 23675 19579 23681
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23681 19671 23715
rect 19613 23675 19671 23681
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23681 19855 23715
rect 19797 23675 19855 23681
rect 16945 23647 17003 23653
rect 16945 23644 16957 23647
rect 16500 23616 16957 23644
rect 16500 23585 16528 23616
rect 16945 23613 16957 23616
rect 16991 23613 17003 23647
rect 16945 23607 17003 23613
rect 18322 23604 18328 23656
rect 18380 23644 18386 23656
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18380 23616 18705 23644
rect 18380 23604 18386 23616
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 18693 23607 18751 23613
rect 16485 23579 16543 23585
rect 16485 23545 16497 23579
rect 16531 23545 16543 23579
rect 16485 23539 16543 23545
rect 16758 23508 16764 23520
rect 16132 23480 16764 23508
rect 14332 23468 14338 23480
rect 16758 23468 16764 23480
rect 16816 23508 16822 23520
rect 18414 23508 18420 23520
rect 16816 23480 18420 23508
rect 16816 23468 16822 23480
rect 18414 23468 18420 23480
rect 18472 23468 18478 23520
rect 18506 23468 18512 23520
rect 18564 23508 18570 23520
rect 18877 23511 18935 23517
rect 18877 23508 18889 23511
rect 18564 23480 18889 23508
rect 18564 23468 18570 23480
rect 18877 23477 18889 23480
rect 18923 23477 18935 23511
rect 18877 23471 18935 23477
rect 19337 23511 19395 23517
rect 19337 23477 19349 23511
rect 19383 23508 19395 23511
rect 19426 23508 19432 23520
rect 19383 23480 19432 23508
rect 19383 23477 19395 23480
rect 19337 23471 19395 23477
rect 19426 23468 19432 23480
rect 19484 23468 19490 23520
rect 19536 23508 19564 23675
rect 19628 23576 19656 23675
rect 19886 23672 19892 23724
rect 19944 23712 19950 23724
rect 20364 23721 20392 23752
rect 22094 23740 22100 23792
rect 22152 23780 22158 23792
rect 23400 23780 23428 23811
rect 23753 23783 23811 23789
rect 23753 23780 23765 23783
rect 22152 23752 23336 23780
rect 23400 23752 23765 23780
rect 22152 23740 22158 23752
rect 20165 23715 20223 23721
rect 20165 23712 20177 23715
rect 19944 23684 20177 23712
rect 19944 23672 19950 23684
rect 20165 23681 20177 23684
rect 20211 23681 20223 23715
rect 20165 23675 20223 23681
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23712 20407 23715
rect 20530 23712 20536 23724
rect 20395 23684 20536 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 22465 23715 22523 23721
rect 22465 23681 22477 23715
rect 22511 23712 22523 23715
rect 22511 23684 23152 23712
rect 22511 23681 22523 23684
rect 22465 23675 22523 23681
rect 20073 23647 20131 23653
rect 20073 23613 20085 23647
rect 20119 23644 20131 23647
rect 20254 23644 20260 23656
rect 20119 23616 20260 23644
rect 20119 23613 20131 23616
rect 20073 23607 20131 23613
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 22370 23604 22376 23656
rect 22428 23604 22434 23656
rect 22830 23604 22836 23656
rect 22888 23604 22894 23656
rect 20898 23576 20904 23588
rect 19628 23548 20904 23576
rect 20898 23536 20904 23548
rect 20956 23536 20962 23588
rect 23124 23576 23152 23684
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 23308 23644 23336 23752
rect 23753 23749 23765 23752
rect 23799 23749 23811 23783
rect 23753 23743 23811 23749
rect 24486 23740 24492 23792
rect 24544 23740 24550 23792
rect 23382 23644 23388 23656
rect 23308 23616 23388 23644
rect 23382 23604 23388 23616
rect 23440 23644 23446 23656
rect 23477 23647 23535 23653
rect 23477 23644 23489 23647
rect 23440 23616 23489 23644
rect 23440 23604 23446 23616
rect 23477 23613 23489 23616
rect 23523 23613 23535 23647
rect 23477 23607 23535 23613
rect 23124 23548 23612 23576
rect 23584 23520 23612 23548
rect 19794 23508 19800 23520
rect 19536 23480 19800 23508
rect 19794 23468 19800 23480
rect 19852 23468 19858 23520
rect 23566 23468 23572 23520
rect 23624 23468 23630 23520
rect 25130 23468 25136 23520
rect 25188 23508 25194 23520
rect 25225 23511 25283 23517
rect 25225 23508 25237 23511
rect 25188 23480 25237 23508
rect 25188 23468 25194 23480
rect 25225 23477 25237 23480
rect 25271 23477 25283 23511
rect 25225 23471 25283 23477
rect 1104 23418 26864 23440
rect 1104 23366 2918 23418
rect 2970 23366 2982 23418
rect 3034 23366 3046 23418
rect 3098 23366 3110 23418
rect 3162 23366 3174 23418
rect 3226 23366 3238 23418
rect 3290 23366 6918 23418
rect 6970 23366 6982 23418
rect 7034 23366 7046 23418
rect 7098 23366 7110 23418
rect 7162 23366 7174 23418
rect 7226 23366 7238 23418
rect 7290 23366 10918 23418
rect 10970 23366 10982 23418
rect 11034 23366 11046 23418
rect 11098 23366 11110 23418
rect 11162 23366 11174 23418
rect 11226 23366 11238 23418
rect 11290 23366 14918 23418
rect 14970 23366 14982 23418
rect 15034 23366 15046 23418
rect 15098 23366 15110 23418
rect 15162 23366 15174 23418
rect 15226 23366 15238 23418
rect 15290 23366 18918 23418
rect 18970 23366 18982 23418
rect 19034 23366 19046 23418
rect 19098 23366 19110 23418
rect 19162 23366 19174 23418
rect 19226 23366 19238 23418
rect 19290 23366 22918 23418
rect 22970 23366 22982 23418
rect 23034 23366 23046 23418
rect 23098 23366 23110 23418
rect 23162 23366 23174 23418
rect 23226 23366 23238 23418
rect 23290 23366 26864 23418
rect 1104 23344 26864 23366
rect 5350 23264 5356 23316
rect 5408 23304 5414 23316
rect 5445 23307 5503 23313
rect 5445 23304 5457 23307
rect 5408 23276 5457 23304
rect 5408 23264 5414 23276
rect 5445 23273 5457 23276
rect 5491 23273 5503 23307
rect 5445 23267 5503 23273
rect 7101 23307 7159 23313
rect 7101 23273 7113 23307
rect 7147 23304 7159 23307
rect 7374 23304 7380 23316
rect 7147 23276 7380 23304
rect 7147 23273 7159 23276
rect 7101 23267 7159 23273
rect 7374 23264 7380 23276
rect 7432 23264 7438 23316
rect 10870 23304 10876 23316
rect 7576 23276 10876 23304
rect 5534 23196 5540 23248
rect 5592 23236 5598 23248
rect 7576 23236 7604 23276
rect 10870 23264 10876 23276
rect 10928 23264 10934 23316
rect 12158 23264 12164 23316
rect 12216 23264 12222 23316
rect 12250 23264 12256 23316
rect 12308 23304 12314 23316
rect 14826 23304 14832 23316
rect 12308 23276 14832 23304
rect 12308 23264 12314 23276
rect 5592 23208 7604 23236
rect 5592 23196 5598 23208
rect 8570 23196 8576 23248
rect 8628 23236 8634 23248
rect 8628 23208 10548 23236
rect 8628 23196 8634 23208
rect 1946 23128 1952 23180
rect 2004 23128 2010 23180
rect 5718 23168 5724 23180
rect 4816 23140 5724 23168
rect 4816 23109 4844 23140
rect 5718 23128 5724 23140
rect 5776 23128 5782 23180
rect 5902 23128 5908 23180
rect 5960 23128 5966 23180
rect 5994 23128 6000 23180
rect 6052 23168 6058 23180
rect 7374 23168 7380 23180
rect 6052 23140 7380 23168
rect 6052 23128 6058 23140
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 8588 23168 8616 23196
rect 8404 23140 8616 23168
rect 4801 23103 4859 23109
rect 4801 23069 4813 23103
rect 4847 23069 4859 23103
rect 4801 23063 4859 23069
rect 5074 23060 5080 23112
rect 5132 23060 5138 23112
rect 5169 23103 5227 23109
rect 5169 23069 5181 23103
rect 5215 23100 5227 23103
rect 5442 23100 5448 23112
rect 5215 23072 5448 23100
rect 5215 23069 5227 23072
rect 5169 23063 5227 23069
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23100 5871 23103
rect 6270 23100 6276 23112
rect 5859 23072 6276 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 6546 23060 6552 23112
rect 6604 23060 6610 23112
rect 6641 23103 6699 23109
rect 6641 23069 6653 23103
rect 6687 23100 6699 23103
rect 8404 23100 8432 23140
rect 9674 23128 9680 23180
rect 9732 23168 9738 23180
rect 10410 23168 10416 23180
rect 9732 23140 10416 23168
rect 9732 23128 9738 23140
rect 10410 23128 10416 23140
rect 10468 23128 10474 23180
rect 10520 23168 10548 23208
rect 12250 23168 12256 23180
rect 10520 23140 12256 23168
rect 12250 23128 12256 23140
rect 12308 23128 12314 23180
rect 6687 23072 8432 23100
rect 8481 23103 8539 23109
rect 6687 23069 6699 23072
rect 6641 23063 6699 23069
rect 8481 23069 8493 23103
rect 8527 23100 8539 23103
rect 8662 23100 8668 23112
rect 8527 23072 8668 23100
rect 8527 23069 8539 23072
rect 8481 23063 8539 23069
rect 8662 23060 8668 23072
rect 8720 23060 8726 23112
rect 8754 23060 8760 23112
rect 8812 23060 8818 23112
rect 9490 23060 9496 23112
rect 9548 23100 9554 23112
rect 9769 23103 9827 23109
rect 9769 23100 9781 23103
rect 9548 23072 9781 23100
rect 9548 23060 9554 23072
rect 9769 23069 9781 23072
rect 9815 23069 9827 23103
rect 9769 23063 9827 23069
rect 10137 23103 10195 23109
rect 10137 23069 10149 23103
rect 10183 23100 10195 23103
rect 10318 23100 10324 23112
rect 10183 23072 10324 23100
rect 10183 23069 10195 23072
rect 10137 23063 10195 23069
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 12360 23100 12388 23276
rect 14826 23264 14832 23276
rect 14884 23304 14890 23316
rect 17310 23304 17316 23316
rect 14884 23276 17316 23304
rect 14884 23264 14890 23276
rect 17310 23264 17316 23276
rect 17368 23264 17374 23316
rect 19886 23304 19892 23316
rect 19260 23276 19892 23304
rect 12434 23196 12440 23248
rect 12492 23236 12498 23248
rect 12492 23208 12572 23236
rect 12492 23196 12498 23208
rect 12544 23177 12572 23208
rect 12529 23171 12587 23177
rect 12529 23137 12541 23171
rect 12575 23137 12587 23171
rect 12529 23131 12587 23137
rect 16666 23128 16672 23180
rect 16724 23128 16730 23180
rect 18414 23128 18420 23180
rect 18472 23168 18478 23180
rect 18693 23171 18751 23177
rect 18693 23168 18705 23171
rect 18472 23140 18705 23168
rect 18472 23128 18478 23140
rect 18693 23137 18705 23140
rect 18739 23137 18751 23171
rect 18693 23131 18751 23137
rect 12437 23103 12495 23109
rect 12437 23100 12449 23103
rect 12360 23072 12449 23100
rect 12437 23069 12449 23072
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12796 23103 12854 23109
rect 12796 23069 12808 23103
rect 12842 23100 12854 23103
rect 13170 23100 13176 23112
rect 12842 23072 13176 23100
rect 12842 23069 12854 23072
rect 12796 23063 12854 23069
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 14090 23060 14096 23112
rect 14148 23060 14154 23112
rect 15562 23060 15568 23112
rect 15620 23100 15626 23112
rect 16114 23109 16120 23112
rect 15933 23103 15991 23109
rect 15933 23100 15945 23103
rect 15620 23072 15945 23100
rect 15620 23060 15626 23072
rect 15933 23069 15945 23072
rect 15979 23069 15991 23103
rect 15933 23063 15991 23069
rect 16081 23103 16120 23109
rect 16081 23069 16093 23103
rect 16081 23063 16120 23069
rect 16114 23060 16120 23063
rect 16172 23060 16178 23112
rect 16298 23060 16304 23112
rect 16356 23060 16362 23112
rect 16439 23103 16497 23109
rect 16439 23069 16451 23103
rect 16485 23100 16497 23103
rect 17402 23100 17408 23112
rect 16485 23072 17408 23100
rect 16485 23069 16497 23072
rect 16439 23063 16497 23069
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 18322 23060 18328 23112
rect 18380 23100 18386 23112
rect 19260 23109 19288 23276
rect 19886 23264 19892 23276
rect 19944 23304 19950 23316
rect 20165 23307 20223 23313
rect 20165 23304 20177 23307
rect 19944 23276 20177 23304
rect 19944 23264 19950 23276
rect 20165 23273 20177 23276
rect 20211 23273 20223 23307
rect 20165 23267 20223 23273
rect 20349 23307 20407 23313
rect 20349 23273 20361 23307
rect 20395 23304 20407 23307
rect 21726 23304 21732 23316
rect 20395 23276 21732 23304
rect 20395 23273 20407 23276
rect 20349 23267 20407 23273
rect 21726 23264 21732 23276
rect 21784 23264 21790 23316
rect 19518 23196 19524 23248
rect 19576 23236 19582 23248
rect 19978 23236 19984 23248
rect 19576 23208 19984 23236
rect 19576 23196 19582 23208
rect 19628 23177 19656 23208
rect 19978 23196 19984 23208
rect 20036 23196 20042 23248
rect 20073 23239 20131 23245
rect 20073 23205 20085 23239
rect 20119 23236 20131 23239
rect 22370 23236 22376 23248
rect 20119 23208 22376 23236
rect 20119 23205 20131 23208
rect 20073 23199 20131 23205
rect 22370 23196 22376 23208
rect 22428 23196 22434 23248
rect 19613 23171 19671 23177
rect 19613 23137 19625 23171
rect 19659 23137 19671 23171
rect 19613 23131 19671 23137
rect 19705 23171 19763 23177
rect 19705 23137 19717 23171
rect 19751 23168 19763 23171
rect 20530 23168 20536 23180
rect 19751 23140 20536 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 20530 23128 20536 23140
rect 20588 23128 20594 23180
rect 22094 23128 22100 23180
rect 22152 23168 22158 23180
rect 22465 23171 22523 23177
rect 22465 23168 22477 23171
rect 22152 23140 22477 23168
rect 22152 23128 22158 23140
rect 22465 23137 22477 23140
rect 22511 23137 22523 23171
rect 22465 23131 22523 23137
rect 22738 23128 22744 23180
rect 22796 23168 22802 23180
rect 22796 23140 24440 23168
rect 22796 23128 22802 23140
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 18380 23072 18521 23100
rect 18380 23060 18386 23072
rect 18509 23069 18521 23072
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 19426 23060 19432 23112
rect 19484 23060 19490 23112
rect 19794 23060 19800 23112
rect 19852 23060 19858 23112
rect 19886 23060 19892 23112
rect 19944 23060 19950 23112
rect 20717 23103 20775 23109
rect 20717 23100 20729 23103
rect 19996 23072 20729 23100
rect 2216 23035 2274 23041
rect 2216 23001 2228 23035
rect 2262 23032 2274 23035
rect 2314 23032 2320 23044
rect 2262 23004 2320 23032
rect 2262 23001 2274 23004
rect 2216 22995 2274 23001
rect 2314 22992 2320 23004
rect 2372 22992 2378 23044
rect 4985 23035 5043 23041
rect 4985 23001 4997 23035
rect 5031 23032 5043 23035
rect 5258 23032 5264 23044
rect 5031 23004 5264 23032
rect 5031 23001 5043 23004
rect 4985 22995 5043 23001
rect 5258 22992 5264 23004
rect 5316 23032 5322 23044
rect 6457 23035 6515 23041
rect 6457 23032 6469 23035
rect 5316 23004 6469 23032
rect 5316 22992 5322 23004
rect 6457 23001 6469 23004
rect 6503 23001 6515 23035
rect 6457 22995 6515 23001
rect 7374 22992 7380 23044
rect 7432 23032 7438 23044
rect 7558 23032 7564 23044
rect 7432 23004 7564 23032
rect 7432 22992 7438 23004
rect 7558 22992 7564 23004
rect 7616 22992 7622 23044
rect 8236 23035 8294 23041
rect 8236 23001 8248 23035
rect 8282 23032 8294 23035
rect 9953 23035 10011 23041
rect 8282 23004 8616 23032
rect 8282 23001 8294 23004
rect 8236 22995 8294 23001
rect 3142 22924 3148 22976
rect 3200 22964 3206 22976
rect 3329 22967 3387 22973
rect 3329 22964 3341 22967
rect 3200 22936 3341 22964
rect 3200 22924 3206 22936
rect 3329 22933 3341 22936
rect 3375 22933 3387 22967
rect 3329 22927 3387 22933
rect 5350 22924 5356 22976
rect 5408 22924 5414 22976
rect 6178 22924 6184 22976
rect 6236 22964 6242 22976
rect 8588 22973 8616 23004
rect 9953 23001 9965 23035
rect 9999 23001 10011 23035
rect 9953 22995 10011 23001
rect 10045 23035 10103 23041
rect 10045 23001 10057 23035
rect 10091 23032 10103 23035
rect 10091 23004 10640 23032
rect 10091 23001 10103 23004
rect 10045 22995 10103 23001
rect 6825 22967 6883 22973
rect 6825 22964 6837 22967
rect 6236 22936 6837 22964
rect 6236 22924 6242 22936
rect 6825 22933 6837 22936
rect 6871 22933 6883 22967
rect 6825 22927 6883 22933
rect 8573 22967 8631 22973
rect 8573 22933 8585 22967
rect 8619 22933 8631 22967
rect 9968 22964 9996 22995
rect 10134 22964 10140 22976
rect 9968 22936 10140 22964
rect 8573 22927 8631 22933
rect 10134 22924 10140 22936
rect 10192 22924 10198 22976
rect 10318 22924 10324 22976
rect 10376 22924 10382 22976
rect 10612 22964 10640 23004
rect 10686 22992 10692 23044
rect 10744 22992 10750 23044
rect 12345 23035 12403 23041
rect 12345 23032 12357 23035
rect 11914 23004 12357 23032
rect 12345 23001 12357 23004
rect 12391 23001 12403 23035
rect 12345 22995 12403 23001
rect 12894 22992 12900 23044
rect 12952 23032 12958 23044
rect 14366 23041 14372 23044
rect 12952 23004 14044 23032
rect 12952 22992 12958 23004
rect 11422 22964 11428 22976
rect 10612 22936 11428 22964
rect 11422 22924 11428 22936
rect 11480 22924 11486 22976
rect 13722 22924 13728 22976
rect 13780 22964 13786 22976
rect 13909 22967 13967 22973
rect 13909 22964 13921 22967
rect 13780 22936 13921 22964
rect 13780 22924 13786 22936
rect 13909 22933 13921 22936
rect 13955 22933 13967 22967
rect 14016 22964 14044 23004
rect 14360 22995 14372 23041
rect 14366 22992 14372 22995
rect 14424 22992 14430 23044
rect 16209 23035 16267 23041
rect 16209 23032 16221 23035
rect 14476 23004 16221 23032
rect 14476 22964 14504 23004
rect 16209 23001 16221 23004
rect 16255 23032 16267 23035
rect 18046 23032 18052 23044
rect 16255 23004 18052 23032
rect 16255 23001 16267 23004
rect 16209 22995 16267 23001
rect 18046 22992 18052 23004
rect 18104 22992 18110 23044
rect 18414 22992 18420 23044
rect 18472 22992 18478 23044
rect 18966 22992 18972 23044
rect 19024 23032 19030 23044
rect 19996 23032 20024 23072
rect 20717 23069 20729 23072
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 20806 23060 20812 23112
rect 20864 23060 20870 23112
rect 20898 23060 20904 23112
rect 20956 23100 20962 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 20956 23072 21189 23100
rect 20956 23060 20962 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 22186 23060 22192 23112
rect 22244 23060 22250 23112
rect 24412 23109 24440 23140
rect 24397 23103 24455 23109
rect 24397 23069 24409 23103
rect 24443 23100 24455 23103
rect 24673 23103 24731 23109
rect 24673 23100 24685 23103
rect 24443 23072 24685 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 24673 23069 24685 23072
rect 24719 23069 24731 23103
rect 24673 23063 24731 23069
rect 19024 23004 20024 23032
rect 20533 23035 20591 23041
rect 19024 22992 19030 23004
rect 20533 23001 20545 23035
rect 20579 23032 20591 23035
rect 21082 23032 21088 23044
rect 20579 23004 21088 23032
rect 20579 23001 20591 23004
rect 20533 22995 20591 23001
rect 21082 22992 21088 23004
rect 21140 22992 21146 23044
rect 22741 23035 22799 23041
rect 22741 23001 22753 23035
rect 22787 23001 22799 23035
rect 24765 23035 24823 23041
rect 24765 23032 24777 23035
rect 23966 23004 24777 23032
rect 22741 22995 22799 23001
rect 24765 23001 24777 23004
rect 24811 23001 24823 23035
rect 24765 22995 24823 23001
rect 14016 22936 14504 22964
rect 13909 22927 13967 22933
rect 15470 22924 15476 22976
rect 15528 22924 15534 22976
rect 16114 22924 16120 22976
rect 16172 22964 16178 22976
rect 16482 22964 16488 22976
rect 16172 22936 16488 22964
rect 16172 22924 16178 22936
rect 16482 22924 16488 22936
rect 16540 22924 16546 22976
rect 16574 22924 16580 22976
rect 16632 22924 16638 22976
rect 19337 22967 19395 22973
rect 19337 22933 19349 22967
rect 19383 22964 19395 22967
rect 19426 22964 19432 22976
rect 19383 22936 19432 22964
rect 19383 22933 19395 22936
rect 19337 22927 19395 22933
rect 19426 22924 19432 22936
rect 19484 22924 19490 22976
rect 20346 22973 20352 22976
rect 20333 22967 20352 22973
rect 20333 22933 20345 22967
rect 20333 22927 20352 22933
rect 20346 22924 20352 22927
rect 20404 22924 20410 22976
rect 20990 22924 20996 22976
rect 21048 22924 21054 22976
rect 22373 22967 22431 22973
rect 22373 22933 22385 22967
rect 22419 22964 22431 22967
rect 22756 22964 22784 22995
rect 22419 22936 22784 22964
rect 22419 22933 22431 22936
rect 22373 22927 22431 22933
rect 24210 22924 24216 22976
rect 24268 22924 24274 22976
rect 24486 22924 24492 22976
rect 24544 22924 24550 22976
rect 1104 22874 26864 22896
rect 1104 22822 3658 22874
rect 3710 22822 3722 22874
rect 3774 22822 3786 22874
rect 3838 22822 3850 22874
rect 3902 22822 3914 22874
rect 3966 22822 3978 22874
rect 4030 22822 7658 22874
rect 7710 22822 7722 22874
rect 7774 22822 7786 22874
rect 7838 22822 7850 22874
rect 7902 22822 7914 22874
rect 7966 22822 7978 22874
rect 8030 22822 11658 22874
rect 11710 22822 11722 22874
rect 11774 22822 11786 22874
rect 11838 22822 11850 22874
rect 11902 22822 11914 22874
rect 11966 22822 11978 22874
rect 12030 22822 15658 22874
rect 15710 22822 15722 22874
rect 15774 22822 15786 22874
rect 15838 22822 15850 22874
rect 15902 22822 15914 22874
rect 15966 22822 15978 22874
rect 16030 22822 19658 22874
rect 19710 22822 19722 22874
rect 19774 22822 19786 22874
rect 19838 22822 19850 22874
rect 19902 22822 19914 22874
rect 19966 22822 19978 22874
rect 20030 22822 23658 22874
rect 23710 22822 23722 22874
rect 23774 22822 23786 22874
rect 23838 22822 23850 22874
rect 23902 22822 23914 22874
rect 23966 22822 23978 22874
rect 24030 22822 26864 22874
rect 1104 22800 26864 22822
rect 2314 22720 2320 22772
rect 2372 22720 2378 22772
rect 2777 22763 2835 22769
rect 2777 22729 2789 22763
rect 2823 22729 2835 22763
rect 2777 22723 2835 22729
rect 2501 22627 2559 22633
rect 2501 22593 2513 22627
rect 2547 22624 2559 22627
rect 2792 22624 2820 22723
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 6549 22763 6607 22769
rect 3200 22732 3740 22760
rect 3200 22720 3206 22732
rect 3237 22695 3295 22701
rect 3237 22661 3249 22695
rect 3283 22692 3295 22695
rect 3326 22692 3332 22704
rect 3283 22664 3332 22692
rect 3283 22661 3295 22664
rect 3237 22655 3295 22661
rect 3326 22652 3332 22664
rect 3384 22652 3390 22704
rect 2547 22596 2820 22624
rect 2547 22593 2559 22596
rect 2501 22587 2559 22593
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 3605 22627 3663 22633
rect 3605 22624 3617 22627
rect 3568 22596 3617 22624
rect 3568 22584 3574 22596
rect 3605 22593 3617 22596
rect 3651 22593 3663 22627
rect 3712 22624 3740 22732
rect 6549 22729 6561 22763
rect 6595 22760 6607 22763
rect 6595 22732 6914 22760
rect 6595 22729 6607 22732
rect 6549 22723 6607 22729
rect 3789 22695 3847 22701
rect 3789 22661 3801 22695
rect 3835 22692 3847 22695
rect 4614 22692 4620 22704
rect 3835 22664 4620 22692
rect 3835 22661 3847 22664
rect 3789 22655 3847 22661
rect 4614 22652 4620 22664
rect 4672 22652 4678 22704
rect 6886 22701 6914 22732
rect 9490 22720 9496 22772
rect 9548 22720 9554 22772
rect 10686 22720 10692 22772
rect 10744 22760 10750 22772
rect 11517 22763 11575 22769
rect 11517 22760 11529 22763
rect 10744 22732 11529 22760
rect 10744 22720 10750 22732
rect 11517 22729 11529 22732
rect 11563 22729 11575 22763
rect 12158 22760 12164 22772
rect 11517 22723 11575 22729
rect 11808 22732 12164 22760
rect 6886 22695 6944 22701
rect 6886 22661 6898 22695
rect 6932 22661 6944 22695
rect 6886 22655 6944 22661
rect 8294 22652 8300 22704
rect 8352 22692 8358 22704
rect 8570 22692 8576 22704
rect 8352 22664 8576 22692
rect 8352 22652 8358 22664
rect 8570 22652 8576 22664
rect 8628 22652 8634 22704
rect 11330 22692 11336 22704
rect 11086 22664 11336 22692
rect 11330 22652 11336 22664
rect 11388 22652 11394 22704
rect 11808 22701 11836 22732
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 13354 22720 13360 22772
rect 13412 22720 13418 22772
rect 13722 22720 13728 22772
rect 13780 22720 13786 22772
rect 14366 22720 14372 22772
rect 14424 22720 14430 22772
rect 14645 22763 14703 22769
rect 14645 22729 14657 22763
rect 14691 22729 14703 22763
rect 14645 22723 14703 22729
rect 15013 22763 15071 22769
rect 15013 22729 15025 22763
rect 15059 22760 15071 22763
rect 15470 22760 15476 22772
rect 15059 22732 15476 22760
rect 15059 22729 15071 22732
rect 15013 22723 15071 22729
rect 11793 22695 11851 22701
rect 11793 22661 11805 22695
rect 11839 22661 11851 22695
rect 11793 22655 11851 22661
rect 12250 22652 12256 22704
rect 12308 22692 12314 22704
rect 12308 22664 12848 22692
rect 12308 22652 12314 22664
rect 3881 22627 3939 22633
rect 3881 22624 3893 22627
rect 3712 22596 3893 22624
rect 3605 22587 3663 22593
rect 3881 22593 3893 22596
rect 3927 22593 3939 22627
rect 3881 22587 3939 22593
rect 3970 22584 3976 22636
rect 4028 22584 4034 22636
rect 6365 22627 6423 22633
rect 6365 22593 6377 22627
rect 6411 22624 6423 22627
rect 7374 22624 7380 22636
rect 6411 22596 7380 22624
rect 6411 22593 6423 22596
rect 6365 22587 6423 22593
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 7466 22584 7472 22636
rect 7524 22624 7530 22636
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7524 22596 8125 22624
rect 7524 22584 7530 22596
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22593 8447 22627
rect 8389 22587 8447 22593
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22624 8539 22627
rect 8754 22624 8760 22636
rect 8527 22596 8760 22624
rect 8527 22593 8539 22596
rect 8481 22587 8539 22593
rect 3421 22559 3479 22565
rect 3421 22525 3433 22559
rect 3467 22556 3479 22559
rect 4430 22556 4436 22568
rect 3467 22528 4436 22556
rect 3467 22525 3479 22528
rect 3421 22519 3479 22525
rect 4430 22516 4436 22528
rect 4488 22516 4494 22568
rect 6454 22516 6460 22568
rect 6512 22556 6518 22568
rect 6641 22559 6699 22565
rect 6641 22556 6653 22559
rect 6512 22528 6653 22556
rect 6512 22516 6518 22528
rect 6641 22525 6653 22528
rect 6687 22525 6699 22559
rect 8404 22556 8432 22587
rect 8754 22584 8760 22596
rect 8812 22584 8818 22636
rect 9309 22627 9367 22633
rect 9309 22624 9321 22627
rect 8956 22596 9321 22624
rect 6641 22519 6699 22525
rect 8036 22528 8432 22556
rect 8036 22432 8064 22528
rect 8956 22488 8984 22596
rect 9309 22593 9321 22596
rect 9355 22593 9367 22627
rect 9309 22587 9367 22593
rect 9582 22584 9588 22636
rect 9640 22584 9646 22636
rect 11701 22627 11759 22633
rect 11701 22624 11713 22627
rect 11072 22596 11713 22624
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22556 9091 22559
rect 9490 22556 9496 22568
rect 9079 22528 9496 22556
rect 9079 22525 9091 22528
rect 9033 22519 9091 22525
rect 9490 22516 9496 22528
rect 9548 22516 9554 22568
rect 9861 22559 9919 22565
rect 9861 22525 9873 22559
rect 9907 22556 9919 22559
rect 10318 22556 10324 22568
rect 9907 22528 10324 22556
rect 9907 22525 9919 22528
rect 9861 22519 9919 22525
rect 10318 22516 10324 22528
rect 10376 22516 10382 22568
rect 10410 22516 10416 22568
rect 10468 22556 10474 22568
rect 11072 22556 11100 22596
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22624 11943 22627
rect 11974 22624 11980 22636
rect 11931 22596 11980 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 11974 22584 11980 22596
rect 12032 22584 12038 22636
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22624 12127 22627
rect 12161 22627 12219 22633
rect 12161 22624 12173 22627
rect 12115 22596 12173 22624
rect 12115 22593 12127 22596
rect 12069 22587 12127 22593
rect 12161 22593 12173 22596
rect 12207 22593 12219 22627
rect 12161 22587 12219 22593
rect 12345 22627 12403 22633
rect 12345 22593 12357 22627
rect 12391 22593 12403 22627
rect 12345 22587 12403 22593
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22593 12771 22627
rect 12713 22587 12771 22593
rect 10468 22528 11100 22556
rect 11333 22559 11391 22565
rect 10468 22516 10474 22528
rect 11333 22525 11345 22559
rect 11379 22556 11391 22559
rect 11422 22556 11428 22568
rect 11379 22528 11428 22556
rect 11379 22525 11391 22528
rect 11333 22519 11391 22525
rect 11422 22516 11428 22528
rect 11480 22516 11486 22568
rect 8956 22460 9260 22488
rect 4157 22423 4215 22429
rect 4157 22389 4169 22423
rect 4203 22420 4215 22423
rect 4522 22420 4528 22432
rect 4203 22392 4528 22420
rect 4203 22389 4215 22392
rect 4157 22383 4215 22389
rect 4522 22380 4528 22392
rect 4580 22380 4586 22432
rect 8018 22380 8024 22432
rect 8076 22380 8082 22432
rect 8665 22423 8723 22429
rect 8665 22389 8677 22423
rect 8711 22420 8723 22423
rect 8846 22420 8852 22432
rect 8711 22392 8852 22420
rect 8711 22389 8723 22392
rect 8665 22383 8723 22389
rect 8846 22380 8852 22392
rect 8904 22380 8910 22432
rect 9122 22380 9128 22432
rect 9180 22380 9186 22432
rect 9232 22420 9260 22460
rect 9950 22420 9956 22432
rect 9232 22392 9956 22420
rect 9950 22380 9956 22392
rect 10008 22420 10014 22432
rect 12360 22420 12388 22587
rect 12618 22516 12624 22568
rect 12676 22516 12682 22568
rect 12728 22488 12756 22587
rect 12820 22556 12848 22664
rect 12894 22652 12900 22704
rect 12952 22652 12958 22704
rect 12989 22695 13047 22701
rect 12989 22661 13001 22695
rect 13035 22692 13047 22695
rect 13740 22692 13768 22720
rect 13035 22664 13768 22692
rect 13035 22661 13047 22664
rect 12989 22655 13047 22661
rect 13081 22627 13139 22633
rect 13081 22593 13093 22627
rect 13127 22593 13139 22627
rect 13081 22587 13139 22593
rect 13096 22556 13124 22587
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 13630 22624 13636 22636
rect 13504 22596 13636 22624
rect 13504 22584 13510 22596
rect 13630 22584 13636 22596
rect 13688 22624 13694 22636
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 13688 22596 13829 22624
rect 13688 22584 13694 22596
rect 13817 22593 13829 22596
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22624 14611 22627
rect 14660 22624 14688 22723
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 20162 22760 20168 22772
rect 16684 22732 20168 22760
rect 16684 22704 16712 22732
rect 15105 22695 15163 22701
rect 15105 22661 15117 22695
rect 15151 22692 15163 22695
rect 16206 22692 16212 22704
rect 15151 22664 16212 22692
rect 15151 22661 15163 22664
rect 15105 22655 15163 22661
rect 16206 22652 16212 22664
rect 16264 22652 16270 22704
rect 16666 22652 16672 22704
rect 16724 22652 16730 22704
rect 17497 22695 17555 22701
rect 17497 22661 17509 22695
rect 17543 22692 17555 22695
rect 17954 22692 17960 22704
rect 17543 22664 17960 22692
rect 17543 22661 17555 22664
rect 17497 22655 17555 22661
rect 17954 22652 17960 22664
rect 18012 22652 18018 22704
rect 18966 22652 18972 22704
rect 19024 22652 19030 22704
rect 19426 22652 19432 22704
rect 19484 22652 19490 22704
rect 16114 22624 16120 22636
rect 14599 22596 14688 22624
rect 14752 22596 16120 22624
rect 14599 22593 14611 22596
rect 14553 22587 14611 22593
rect 12820 22528 13124 22556
rect 13538 22516 13544 22568
rect 13596 22556 13602 22568
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 13596 22528 14013 22556
rect 13596 22516 13602 22528
rect 14001 22525 14013 22528
rect 14047 22556 14059 22559
rect 14752 22556 14780 22596
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 17310 22584 17316 22636
rect 17368 22624 17374 22636
rect 19720 22633 19748 22732
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 22186 22720 22192 22772
rect 22244 22760 22250 22772
rect 22741 22763 22799 22769
rect 22741 22760 22753 22763
rect 22244 22732 22753 22760
rect 22244 22720 22250 22732
rect 22741 22729 22753 22732
rect 22787 22729 22799 22763
rect 22741 22723 22799 22729
rect 20070 22652 20076 22704
rect 20128 22692 20134 22704
rect 22373 22695 22431 22701
rect 20128 22664 20300 22692
rect 20128 22652 20134 22664
rect 17405 22627 17463 22633
rect 17405 22624 17417 22627
rect 17368 22596 17417 22624
rect 17368 22584 17374 22596
rect 17405 22593 17417 22596
rect 17451 22593 17463 22627
rect 17405 22587 17463 22593
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22593 19763 22627
rect 20162 22624 20168 22636
rect 19705 22587 19763 22593
rect 20088 22596 20168 22624
rect 14047 22528 14780 22556
rect 15197 22559 15255 22565
rect 14047 22525 14059 22528
rect 14001 22519 14059 22525
rect 15197 22525 15209 22559
rect 15243 22525 15255 22559
rect 15197 22519 15255 22525
rect 14274 22488 14280 22500
rect 12728 22460 14280 22488
rect 14274 22448 14280 22460
rect 14332 22448 14338 22500
rect 14826 22448 14832 22500
rect 14884 22488 14890 22500
rect 15212 22488 15240 22519
rect 14884 22460 15240 22488
rect 14884 22448 14890 22460
rect 10008 22392 12388 22420
rect 12529 22423 12587 22429
rect 10008 22380 10014 22392
rect 12529 22389 12541 22423
rect 12575 22420 12587 22423
rect 12710 22420 12716 22432
rect 12575 22392 12716 22420
rect 12575 22389 12587 22392
rect 12529 22383 12587 22389
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 13265 22423 13323 22429
rect 13265 22389 13277 22423
rect 13311 22420 13323 22423
rect 13722 22420 13728 22432
rect 13311 22392 13728 22420
rect 13311 22389 13323 22392
rect 13265 22383 13323 22389
rect 13722 22380 13728 22392
rect 13780 22380 13786 22432
rect 17420 22420 17448 22587
rect 17678 22516 17684 22568
rect 17736 22516 17742 22568
rect 20088 22565 20116 22596
rect 20162 22584 20168 22596
rect 20220 22584 20226 22636
rect 20272 22633 20300 22664
rect 22373 22661 22385 22695
rect 22419 22692 22431 22695
rect 24210 22692 24216 22704
rect 22419 22664 24216 22692
rect 22419 22661 22431 22664
rect 22373 22655 22431 22661
rect 24210 22652 24216 22664
rect 24268 22652 24274 22704
rect 24486 22652 24492 22704
rect 24544 22652 24550 22704
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22593 20315 22627
rect 20257 22587 20315 22593
rect 20438 22584 20444 22636
rect 20496 22624 20502 22636
rect 20533 22627 20591 22633
rect 20533 22624 20545 22627
rect 20496 22596 20545 22624
rect 20496 22584 20502 22596
rect 20533 22593 20545 22596
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 20809 22627 20867 22633
rect 20809 22593 20821 22627
rect 20855 22624 20867 22627
rect 21082 22624 21088 22636
rect 20855 22596 21088 22624
rect 20855 22593 20867 22596
rect 20809 22587 20867 22593
rect 21082 22584 21088 22596
rect 21140 22584 21146 22636
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22624 21419 22627
rect 21726 22624 21732 22636
rect 21407 22596 21732 22624
rect 21407 22593 21419 22596
rect 21361 22587 21419 22593
rect 21726 22584 21732 22596
rect 21784 22584 21790 22636
rect 23382 22584 23388 22636
rect 23440 22624 23446 22636
rect 23661 22627 23719 22633
rect 23661 22624 23673 22627
rect 23440 22596 23673 22624
rect 23440 22584 23446 22596
rect 23661 22593 23673 22596
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 25222 22584 25228 22636
rect 25280 22624 25286 22636
rect 26329 22627 26387 22633
rect 26329 22624 26341 22627
rect 25280 22596 26341 22624
rect 25280 22584 25286 22596
rect 26329 22593 26341 22596
rect 26375 22593 26387 22627
rect 26329 22587 26387 22593
rect 20073 22559 20131 22565
rect 20073 22525 20085 22559
rect 20119 22525 20131 22559
rect 20714 22556 20720 22568
rect 20073 22519 20131 22525
rect 20272 22528 20720 22556
rect 20272 22420 20300 22528
rect 20714 22516 20720 22528
rect 20772 22516 20778 22568
rect 21100 22556 21128 22584
rect 21542 22556 21548 22568
rect 21100 22528 21548 22556
rect 21542 22516 21548 22528
rect 21600 22516 21606 22568
rect 22189 22559 22247 22565
rect 22189 22525 22201 22559
rect 22235 22525 22247 22559
rect 22189 22519 22247 22525
rect 20441 22491 20499 22497
rect 20441 22457 20453 22491
rect 20487 22488 20499 22491
rect 20530 22488 20536 22500
rect 20487 22460 20536 22488
rect 20487 22457 20499 22460
rect 20441 22451 20499 22457
rect 17420 22392 20300 22420
rect 20346 22380 20352 22432
rect 20404 22420 20410 22432
rect 20456 22420 20484 22451
rect 20530 22448 20536 22460
rect 20588 22448 20594 22500
rect 21174 22448 21180 22500
rect 21232 22488 21238 22500
rect 21269 22491 21327 22497
rect 21269 22488 21281 22491
rect 21232 22460 21281 22488
rect 21232 22448 21238 22460
rect 21269 22457 21281 22460
rect 21315 22457 21327 22491
rect 21269 22451 21327 22457
rect 21910 22448 21916 22500
rect 21968 22488 21974 22500
rect 22204 22488 22232 22519
rect 22278 22516 22284 22568
rect 22336 22516 22342 22568
rect 23934 22516 23940 22568
rect 23992 22516 23998 22568
rect 23474 22488 23480 22500
rect 21968 22460 23480 22488
rect 21968 22448 21974 22460
rect 23474 22448 23480 22460
rect 23532 22448 23538 22500
rect 26510 22448 26516 22500
rect 26568 22448 26574 22500
rect 20404 22392 20484 22420
rect 20404 22380 20410 22392
rect 25406 22380 25412 22432
rect 25464 22380 25470 22432
rect 1104 22330 26864 22352
rect 1104 22278 2918 22330
rect 2970 22278 2982 22330
rect 3034 22278 3046 22330
rect 3098 22278 3110 22330
rect 3162 22278 3174 22330
rect 3226 22278 3238 22330
rect 3290 22278 6918 22330
rect 6970 22278 6982 22330
rect 7034 22278 7046 22330
rect 7098 22278 7110 22330
rect 7162 22278 7174 22330
rect 7226 22278 7238 22330
rect 7290 22278 10918 22330
rect 10970 22278 10982 22330
rect 11034 22278 11046 22330
rect 11098 22278 11110 22330
rect 11162 22278 11174 22330
rect 11226 22278 11238 22330
rect 11290 22278 14918 22330
rect 14970 22278 14982 22330
rect 15034 22278 15046 22330
rect 15098 22278 15110 22330
rect 15162 22278 15174 22330
rect 15226 22278 15238 22330
rect 15290 22278 18918 22330
rect 18970 22278 18982 22330
rect 19034 22278 19046 22330
rect 19098 22278 19110 22330
rect 19162 22278 19174 22330
rect 19226 22278 19238 22330
rect 19290 22278 22918 22330
rect 22970 22278 22982 22330
rect 23034 22278 23046 22330
rect 23098 22278 23110 22330
rect 23162 22278 23174 22330
rect 23226 22278 23238 22330
rect 23290 22278 26864 22330
rect 1104 22256 26864 22278
rect 7193 22219 7251 22225
rect 7193 22185 7205 22219
rect 7239 22216 7251 22219
rect 7374 22216 7380 22228
rect 7239 22188 7380 22216
rect 7239 22185 7251 22188
rect 7193 22179 7251 22185
rect 7374 22176 7380 22188
rect 7432 22176 7438 22228
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 12437 22219 12495 22225
rect 9180 22188 12020 22216
rect 9180 22176 9186 22188
rect 3970 22108 3976 22160
rect 4028 22148 4034 22160
rect 4246 22148 4252 22160
rect 4028 22120 4252 22148
rect 4028 22108 4034 22120
rect 4246 22108 4252 22120
rect 4304 22148 4310 22160
rect 8754 22148 8760 22160
rect 4304 22120 8760 22148
rect 4304 22108 4310 22120
rect 8754 22108 8760 22120
rect 8812 22108 8818 22160
rect 11992 22148 12020 22188
rect 12437 22185 12449 22219
rect 12483 22216 12495 22219
rect 12618 22216 12624 22228
rect 12483 22188 12624 22216
rect 12483 22185 12495 22188
rect 12437 22179 12495 22185
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 15749 22219 15807 22225
rect 15749 22216 15761 22219
rect 15620 22188 15761 22216
rect 15620 22176 15626 22188
rect 15749 22185 15761 22188
rect 15795 22185 15807 22219
rect 15749 22179 15807 22185
rect 17862 22176 17868 22228
rect 17920 22216 17926 22228
rect 19518 22216 19524 22228
rect 17920 22188 19524 22216
rect 17920 22176 17926 22188
rect 19518 22176 19524 22188
rect 19576 22176 19582 22228
rect 20070 22176 20076 22228
rect 20128 22216 20134 22228
rect 21361 22219 21419 22225
rect 20128 22188 20760 22216
rect 20128 22176 20134 22188
rect 12710 22148 12716 22160
rect 11992 22120 12716 22148
rect 12710 22108 12716 22120
rect 12768 22148 12774 22160
rect 13906 22148 13912 22160
rect 12768 22120 13912 22148
rect 12768 22108 12774 22120
rect 13906 22108 13912 22120
rect 13964 22108 13970 22160
rect 18616 22120 20668 22148
rect 4338 22040 4344 22092
rect 4396 22080 4402 22092
rect 6454 22080 6460 22092
rect 4396 22052 6460 22080
rect 4396 22040 4402 22052
rect 6454 22040 6460 22052
rect 6512 22040 6518 22092
rect 7837 22083 7895 22089
rect 7837 22049 7849 22083
rect 7883 22080 7895 22083
rect 8202 22080 8208 22092
rect 7883 22052 8208 22080
rect 7883 22049 7895 22052
rect 7837 22043 7895 22049
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 8662 22040 8668 22092
rect 8720 22080 8726 22092
rect 8941 22083 8999 22089
rect 8941 22080 8953 22083
rect 8720 22052 8953 22080
rect 8720 22040 8726 22052
rect 8941 22049 8953 22052
rect 8987 22049 8999 22083
rect 8941 22043 8999 22049
rect 2682 21972 2688 22024
rect 2740 21972 2746 22024
rect 4890 21972 4896 22024
rect 4948 21972 4954 22024
rect 5166 21972 5172 22024
rect 5224 21972 5230 22024
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 22012 5411 22015
rect 7561 22015 7619 22021
rect 5399 21984 5433 22012
rect 5399 21981 5411 21984
rect 5353 21975 5411 21981
rect 7561 21981 7573 22015
rect 7607 22012 7619 22015
rect 8018 22012 8024 22024
rect 7607 21984 8024 22012
rect 7607 21981 7619 21984
rect 7561 21975 7619 21981
rect 4614 21904 4620 21956
rect 4672 21944 4678 21956
rect 5368 21944 5396 21975
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 8570 21972 8576 22024
rect 8628 21972 8634 22024
rect 8956 22012 8984 22043
rect 15470 22040 15476 22092
rect 15528 22040 15534 22092
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 17368 22052 18153 22080
rect 17368 22040 17374 22052
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 18141 22043 18199 22049
rect 11057 22015 11115 22021
rect 11057 22012 11069 22015
rect 8956 21984 11069 22012
rect 11057 21981 11069 21984
rect 11103 22012 11115 22015
rect 12434 22012 12440 22024
rect 11103 21984 12440 22012
rect 11103 21981 11115 21984
rect 11057 21975 11115 21981
rect 12434 21972 12440 21984
rect 12492 21972 12498 22024
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 22012 15255 22015
rect 15488 22012 15516 22040
rect 15243 21984 15516 22012
rect 15243 21981 15255 21984
rect 15197 21975 15255 21981
rect 15562 21972 15568 22024
rect 15620 21972 15626 22024
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 5442 21944 5448 21956
rect 4672 21916 5448 21944
rect 4672 21904 4678 21916
rect 5442 21904 5448 21916
rect 5500 21904 5506 21956
rect 9186 21947 9244 21953
rect 9186 21944 9198 21947
rect 8772 21916 9198 21944
rect 2314 21836 2320 21888
rect 2372 21876 2378 21888
rect 2501 21879 2559 21885
rect 2501 21876 2513 21879
rect 2372 21848 2513 21876
rect 2372 21836 2378 21848
rect 2501 21845 2513 21848
rect 2547 21845 2559 21879
rect 2501 21839 2559 21845
rect 4706 21836 4712 21888
rect 4764 21836 4770 21888
rect 5537 21879 5595 21885
rect 5537 21845 5549 21879
rect 5583 21876 5595 21879
rect 5902 21876 5908 21888
rect 5583 21848 5908 21876
rect 5583 21845 5595 21848
rect 5537 21839 5595 21845
rect 5902 21836 5908 21848
rect 5960 21836 5966 21888
rect 7653 21879 7711 21885
rect 7653 21845 7665 21879
rect 7699 21876 7711 21879
rect 8110 21876 8116 21888
rect 7699 21848 8116 21876
rect 7699 21845 7711 21848
rect 7653 21839 7711 21845
rect 8110 21836 8116 21848
rect 8168 21836 8174 21888
rect 8772 21885 8800 21916
rect 9186 21913 9198 21916
rect 9232 21913 9244 21947
rect 9186 21907 9244 21913
rect 11146 21904 11152 21956
rect 11204 21944 11210 21956
rect 11302 21947 11360 21953
rect 11302 21944 11314 21947
rect 11204 21916 11314 21944
rect 11204 21904 11210 21916
rect 11302 21913 11314 21916
rect 11348 21913 11360 21947
rect 11302 21907 11360 21913
rect 15378 21904 15384 21956
rect 15436 21904 15442 21956
rect 15470 21904 15476 21956
rect 15528 21904 15534 21956
rect 16316 21944 16344 21975
rect 16758 21972 16764 22024
rect 16816 22012 16822 22024
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16816 21984 16865 22012
rect 16816 21972 16822 21984
rect 16853 21981 16865 21984
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 17773 22015 17831 22021
rect 17773 21981 17785 22015
rect 17819 22012 17831 22015
rect 18506 22012 18512 22024
rect 17819 21984 18512 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 17126 21944 17132 21956
rect 16316 21916 17132 21944
rect 17126 21904 17132 21916
rect 17184 21904 17190 21956
rect 17420 21944 17448 21975
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 17586 21944 17592 21956
rect 17420 21916 17592 21944
rect 17586 21904 17592 21916
rect 17644 21944 17650 21956
rect 17862 21944 17868 21956
rect 17644 21916 17868 21944
rect 17644 21904 17650 21916
rect 17862 21904 17868 21916
rect 17920 21944 17926 21956
rect 18049 21947 18107 21953
rect 18049 21944 18061 21947
rect 17920 21916 18061 21944
rect 17920 21904 17926 21916
rect 18049 21913 18061 21916
rect 18095 21913 18107 21947
rect 18049 21907 18107 21913
rect 18322 21904 18328 21956
rect 18380 21944 18386 21956
rect 18616 21953 18644 22120
rect 19242 22040 19248 22092
rect 19300 22080 19306 22092
rect 19300 22052 20024 22080
rect 19300 22040 19306 22052
rect 18690 21972 18696 22024
rect 18748 22012 18754 22024
rect 19061 22015 19119 22021
rect 19061 22012 19073 22015
rect 18748 21984 19073 22012
rect 18748 21972 18754 21984
rect 19061 21981 19073 21984
rect 19107 22012 19119 22015
rect 19797 22015 19855 22021
rect 19352 22012 19564 22014
rect 19797 22012 19809 22015
rect 19107 21986 19809 22012
rect 19107 21984 19380 21986
rect 19536 21984 19809 21986
rect 19107 21981 19119 21984
rect 19061 21975 19119 21981
rect 19797 21981 19809 21984
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 19886 21972 19892 22024
rect 19944 21972 19950 22024
rect 18601 21947 18659 21953
rect 18601 21944 18613 21947
rect 18380 21916 18613 21944
rect 18380 21904 18386 21916
rect 18601 21913 18613 21916
rect 18647 21913 18659 21947
rect 19337 21947 19395 21953
rect 19337 21944 19349 21947
rect 18601 21907 18659 21913
rect 19260 21916 19349 21944
rect 8757 21879 8815 21885
rect 8757 21845 8769 21879
rect 8803 21845 8815 21879
rect 8757 21839 8815 21845
rect 9490 21836 9496 21888
rect 9548 21876 9554 21888
rect 10321 21879 10379 21885
rect 10321 21876 10333 21879
rect 9548 21848 10333 21876
rect 9548 21836 9554 21848
rect 10321 21845 10333 21848
rect 10367 21845 10379 21879
rect 15396 21876 15424 21904
rect 16485 21879 16543 21885
rect 16485 21876 16497 21879
rect 15396 21848 16497 21876
rect 10321 21839 10379 21845
rect 16485 21845 16497 21848
rect 16531 21845 16543 21879
rect 16485 21839 16543 21845
rect 17678 21836 17684 21888
rect 17736 21876 17742 21888
rect 19260 21876 19288 21916
rect 19337 21913 19349 21916
rect 19383 21913 19395 21947
rect 19337 21907 19395 21913
rect 19429 21947 19487 21953
rect 19429 21913 19441 21947
rect 19475 21944 19487 21947
rect 19996 21944 20024 22052
rect 20070 21972 20076 22024
rect 20128 22012 20134 22024
rect 20640 22021 20668 22120
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 20128 21984 20361 22012
rect 20128 21972 20134 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 21981 20591 22015
rect 20533 21975 20591 21981
rect 20625 22015 20683 22021
rect 20625 21981 20637 22015
rect 20671 21981 20683 22015
rect 20732 22012 20760 22188
rect 21361 22185 21373 22219
rect 21407 22216 21419 22219
rect 22278 22216 22284 22228
rect 21407 22188 22284 22216
rect 21407 22185 21419 22188
rect 21361 22179 21419 22185
rect 22278 22176 22284 22188
rect 22336 22176 22342 22228
rect 23934 22176 23940 22228
rect 23992 22216 23998 22228
rect 24029 22219 24087 22225
rect 24029 22216 24041 22219
rect 23992 22188 24041 22216
rect 23992 22176 23998 22188
rect 24029 22185 24041 22188
rect 24075 22185 24087 22219
rect 24029 22179 24087 22185
rect 20898 22108 20904 22160
rect 20956 22148 20962 22160
rect 21910 22148 21916 22160
rect 20956 22120 21916 22148
rect 20956 22108 20962 22120
rect 21910 22108 21916 22120
rect 21968 22108 21974 22160
rect 23474 22148 23480 22160
rect 23400 22120 23480 22148
rect 23400 22089 23428 22120
rect 23474 22108 23480 22120
rect 23532 22108 23538 22160
rect 21177 22083 21235 22089
rect 21177 22049 21189 22083
rect 21223 22080 21235 22083
rect 22097 22083 22155 22089
rect 22097 22080 22109 22083
rect 21223 22052 22109 22080
rect 21223 22049 21235 22052
rect 21177 22043 21235 22049
rect 22097 22049 22109 22052
rect 22143 22049 22155 22083
rect 22097 22043 22155 22049
rect 23385 22083 23443 22089
rect 23385 22049 23397 22083
rect 23431 22080 23443 22083
rect 24489 22083 24547 22089
rect 23431 22052 23465 22080
rect 23431 22049 23443 22052
rect 23385 22043 23443 22049
rect 24489 22049 24501 22083
rect 24535 22080 24547 22083
rect 25222 22080 25228 22092
rect 24535 22052 25228 22080
rect 24535 22049 24547 22052
rect 24489 22043 24547 22049
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 21085 22015 21143 22021
rect 21085 22012 21097 22015
rect 20732 21984 21097 22012
rect 20625 21975 20683 21981
rect 21085 21981 21097 21984
rect 21131 21981 21143 22015
rect 21085 21975 21143 21981
rect 19475 21916 20024 21944
rect 19475 21913 19487 21916
rect 19429 21907 19487 21913
rect 19518 21876 19524 21888
rect 17736 21848 19524 21876
rect 17736 21836 17742 21848
rect 19518 21836 19524 21848
rect 19576 21876 19582 21888
rect 20548 21876 20576 21975
rect 21542 21972 21548 22024
rect 21600 21972 21606 22024
rect 21726 21972 21732 22024
rect 21784 21972 21790 22024
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22020 21944 22048 21975
rect 22186 21972 22192 22024
rect 22244 21972 22250 22024
rect 24213 22015 24271 22021
rect 24213 21981 24225 22015
rect 24259 21981 24271 22015
rect 24213 21975 24271 21981
rect 20824 21916 22048 21944
rect 23569 21947 23627 21953
rect 20824 21888 20852 21916
rect 23569 21913 23581 21947
rect 23615 21944 23627 21947
rect 24118 21944 24124 21956
rect 23615 21916 24124 21944
rect 23615 21913 23627 21916
rect 23569 21907 23627 21913
rect 24118 21904 24124 21916
rect 24176 21904 24182 21956
rect 19576 21848 20576 21876
rect 19576 21836 19582 21848
rect 20806 21836 20812 21888
rect 20864 21836 20870 21888
rect 23474 21836 23480 21888
rect 23532 21836 23538 21888
rect 23937 21879 23995 21885
rect 23937 21845 23949 21879
rect 23983 21876 23995 21879
rect 24228 21876 24256 21975
rect 24394 21972 24400 22024
rect 24452 21972 24458 22024
rect 23983 21848 24256 21876
rect 23983 21845 23995 21848
rect 23937 21839 23995 21845
rect 1104 21786 26864 21808
rect 1104 21734 3658 21786
rect 3710 21734 3722 21786
rect 3774 21734 3786 21786
rect 3838 21734 3850 21786
rect 3902 21734 3914 21786
rect 3966 21734 3978 21786
rect 4030 21734 7658 21786
rect 7710 21734 7722 21786
rect 7774 21734 7786 21786
rect 7838 21734 7850 21786
rect 7902 21734 7914 21786
rect 7966 21734 7978 21786
rect 8030 21734 11658 21786
rect 11710 21734 11722 21786
rect 11774 21734 11786 21786
rect 11838 21734 11850 21786
rect 11902 21734 11914 21786
rect 11966 21734 11978 21786
rect 12030 21734 15658 21786
rect 15710 21734 15722 21786
rect 15774 21734 15786 21786
rect 15838 21734 15850 21786
rect 15902 21734 15914 21786
rect 15966 21734 15978 21786
rect 16030 21734 19658 21786
rect 19710 21734 19722 21786
rect 19774 21734 19786 21786
rect 19838 21734 19850 21786
rect 19902 21734 19914 21786
rect 19966 21734 19978 21786
rect 20030 21734 23658 21786
rect 23710 21734 23722 21786
rect 23774 21734 23786 21786
rect 23838 21734 23850 21786
rect 23902 21734 23914 21786
rect 23966 21734 23978 21786
rect 24030 21734 26864 21786
rect 1104 21712 26864 21734
rect 7009 21675 7067 21681
rect 7009 21672 7021 21675
rect 6196 21644 7021 21672
rect 4516 21607 4574 21613
rect 2056 21576 2774 21604
rect 1946 21496 1952 21548
rect 2004 21536 2010 21548
rect 2056 21545 2084 21576
rect 2314 21545 2320 21548
rect 2041 21539 2099 21545
rect 2041 21536 2053 21539
rect 2004 21508 2053 21536
rect 2004 21496 2010 21508
rect 2041 21505 2053 21508
rect 2087 21505 2099 21539
rect 2308 21536 2320 21545
rect 2275 21508 2320 21536
rect 2041 21499 2099 21505
rect 2308 21499 2320 21508
rect 2314 21496 2320 21499
rect 2372 21496 2378 21548
rect 2746 21536 2774 21576
rect 4516 21573 4528 21607
rect 4562 21604 4574 21607
rect 4706 21604 4712 21616
rect 4562 21576 4712 21604
rect 4562 21573 4574 21576
rect 4516 21567 4574 21573
rect 4706 21564 4712 21576
rect 4764 21564 4770 21616
rect 5350 21564 5356 21616
rect 5408 21604 5414 21616
rect 6196 21613 6224 21644
rect 7009 21641 7021 21644
rect 7055 21641 7067 21675
rect 7009 21635 7067 21641
rect 8570 21632 8576 21684
rect 8628 21672 8634 21684
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 8628 21644 9137 21672
rect 8628 21632 8634 21644
rect 9125 21641 9137 21644
rect 9171 21641 9183 21675
rect 9125 21635 9183 21641
rect 9490 21632 9496 21684
rect 9548 21632 9554 21684
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 11517 21675 11575 21681
rect 11517 21641 11529 21675
rect 11563 21641 11575 21675
rect 11517 21635 11575 21641
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12618 21672 12624 21684
rect 11931 21644 12624 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 6181 21607 6239 21613
rect 5408 21576 6040 21604
rect 5408 21564 5414 21576
rect 4249 21539 4307 21545
rect 4249 21536 4261 21539
rect 2746 21508 4261 21536
rect 4249 21505 4261 21508
rect 4295 21536 4307 21539
rect 4338 21536 4344 21548
rect 4295 21508 4344 21536
rect 4295 21505 4307 21508
rect 4249 21499 4307 21505
rect 4338 21496 4344 21508
rect 4396 21496 4402 21548
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 6012 21536 6040 21576
rect 6181 21573 6193 21607
rect 6227 21573 6239 21607
rect 6733 21607 6791 21613
rect 6733 21604 6745 21607
rect 6181 21567 6239 21573
rect 6279 21576 6745 21604
rect 6279 21536 6307 21576
rect 6733 21573 6745 21576
rect 6779 21573 6791 21607
rect 6733 21567 6791 21573
rect 8202 21564 8208 21616
rect 8260 21604 8266 21616
rect 10042 21604 10048 21616
rect 8260 21576 10048 21604
rect 8260 21564 8266 21576
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 6012 21508 6307 21536
rect 6362 21496 6368 21548
rect 6420 21496 6426 21548
rect 6458 21539 6516 21545
rect 6458 21505 6470 21539
rect 6504 21505 6516 21539
rect 6458 21499 6516 21505
rect 5994 21428 6000 21480
rect 6052 21428 6058 21480
rect 6472 21400 6500 21499
rect 6638 21496 6644 21548
rect 6696 21496 6702 21548
rect 6822 21496 6828 21548
rect 6880 21545 6886 21548
rect 6880 21499 6888 21545
rect 6880 21496 6886 21499
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 11333 21539 11391 21545
rect 8996 21508 9720 21536
rect 8996 21496 9002 21508
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 9692 21477 9720 21508
rect 11333 21505 11345 21539
rect 11379 21536 11391 21539
rect 11532 21536 11560 21635
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 15470 21632 15476 21684
rect 15528 21672 15534 21684
rect 15565 21675 15623 21681
rect 15565 21672 15577 21675
rect 15528 21644 15577 21672
rect 15528 21632 15534 21644
rect 15565 21641 15577 21644
rect 15611 21672 15623 21675
rect 16025 21675 16083 21681
rect 16025 21672 16037 21675
rect 15611 21644 16037 21672
rect 15611 21641 15623 21644
rect 15565 21635 15623 21641
rect 16025 21641 16037 21644
rect 16071 21641 16083 21675
rect 16025 21635 16083 21641
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 19242 21672 19248 21684
rect 18012 21644 19248 21672
rect 18012 21632 18018 21644
rect 19242 21632 19248 21644
rect 19300 21632 19306 21684
rect 19610 21632 19616 21684
rect 19668 21672 19674 21684
rect 21266 21672 21272 21684
rect 19668 21644 21272 21672
rect 19668 21632 19674 21644
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 21726 21632 21732 21684
rect 21784 21672 21790 21684
rect 24394 21672 24400 21684
rect 21784 21644 24400 21672
rect 21784 21632 21790 21644
rect 24394 21632 24400 21644
rect 24452 21632 24458 21684
rect 19797 21607 19855 21613
rect 19797 21573 19809 21607
rect 19843 21604 19855 21607
rect 20530 21604 20536 21616
rect 19843 21576 20536 21604
rect 19843 21573 19855 21576
rect 19797 21567 19855 21573
rect 20530 21564 20536 21576
rect 20588 21564 20594 21616
rect 22186 21604 22192 21616
rect 20640 21576 22192 21604
rect 11379 21508 11560 21536
rect 11977 21539 12035 21545
rect 11379 21505 11391 21508
rect 11333 21499 11391 21505
rect 11977 21505 11989 21539
rect 12023 21536 12035 21539
rect 12250 21536 12256 21548
rect 12023 21508 12256 21536
rect 12023 21505 12035 21508
rect 11977 21499 12035 21505
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 14090 21496 14096 21548
rect 14148 21536 14154 21548
rect 14458 21545 14464 21548
rect 14185 21539 14243 21545
rect 14185 21536 14197 21539
rect 14148 21508 14197 21536
rect 14148 21496 14154 21508
rect 14185 21505 14197 21508
rect 14231 21505 14243 21539
rect 14185 21499 14243 21505
rect 14452 21499 14464 21545
rect 14458 21496 14464 21499
rect 14516 21496 14522 21548
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 16298 21536 16304 21548
rect 16163 21508 16304 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 16298 21496 16304 21508
rect 16356 21496 16362 21548
rect 19981 21539 20039 21545
rect 19981 21505 19993 21539
rect 20027 21505 20039 21539
rect 19981 21499 20039 21505
rect 9585 21471 9643 21477
rect 9585 21468 9597 21471
rect 9456 21440 9597 21468
rect 9456 21428 9462 21440
rect 9585 21437 9597 21440
rect 9631 21437 9643 21471
rect 9585 21431 9643 21437
rect 9677 21471 9735 21477
rect 9677 21437 9689 21471
rect 9723 21437 9735 21471
rect 9677 21431 9735 21437
rect 12069 21471 12127 21477
rect 12069 21437 12081 21471
rect 12115 21468 12127 21471
rect 12342 21468 12348 21480
rect 12115 21440 12348 21468
rect 12115 21437 12127 21440
rect 12069 21431 12127 21437
rect 5644 21372 6500 21400
rect 9692 21400 9720 21431
rect 12084 21400 12112 21431
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 16206 21428 16212 21480
rect 16264 21428 16270 21480
rect 18598 21428 18604 21480
rect 18656 21468 18662 21480
rect 19996 21468 20024 21499
rect 20346 21496 20352 21548
rect 20404 21536 20410 21548
rect 20640 21545 20668 21576
rect 22186 21564 22192 21576
rect 22244 21564 22250 21616
rect 20625 21539 20683 21545
rect 20625 21536 20637 21539
rect 20404 21508 20637 21536
rect 20404 21496 20410 21508
rect 20625 21505 20637 21508
rect 20671 21505 20683 21539
rect 20625 21499 20683 21505
rect 21174 21496 21180 21548
rect 21232 21496 21238 21548
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21536 22063 21539
rect 22646 21536 22652 21548
rect 22051 21508 22652 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24762 21536 24768 21548
rect 24351 21508 24768 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 25133 21539 25191 21545
rect 25133 21505 25145 21539
rect 25179 21536 25191 21539
rect 25406 21536 25412 21548
rect 25179 21508 25412 21536
rect 25179 21505 25191 21508
rect 25133 21499 25191 21505
rect 18656 21440 20376 21468
rect 18656 21428 18662 21440
rect 9692 21372 12112 21400
rect 5644 21344 5672 21372
rect 18414 21360 18420 21412
rect 18472 21400 18478 21412
rect 18509 21403 18567 21409
rect 18509 21400 18521 21403
rect 18472 21372 18521 21400
rect 18472 21360 18478 21372
rect 18509 21369 18521 21372
rect 18555 21400 18567 21403
rect 20254 21400 20260 21412
rect 18555 21372 20260 21400
rect 18555 21369 18567 21372
rect 18509 21363 18567 21369
rect 20254 21360 20260 21372
rect 20312 21360 20318 21412
rect 20348 21400 20376 21440
rect 20530 21428 20536 21480
rect 20588 21428 20594 21480
rect 20993 21471 21051 21477
rect 20993 21437 21005 21471
rect 21039 21468 21051 21471
rect 23474 21468 23480 21480
rect 21039 21440 23480 21468
rect 21039 21437 21051 21440
rect 20993 21431 21051 21437
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 24118 21428 24124 21480
rect 24176 21468 24182 21480
rect 24578 21468 24584 21480
rect 24176 21440 24584 21468
rect 24176 21428 24182 21440
rect 24578 21428 24584 21440
rect 24636 21468 24642 21480
rect 25148 21468 25176 21499
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 25777 21539 25835 21545
rect 25777 21505 25789 21539
rect 25823 21536 25835 21539
rect 26050 21536 26056 21548
rect 25823 21508 26056 21536
rect 25823 21505 25835 21508
rect 25777 21499 25835 21505
rect 26050 21496 26056 21508
rect 26108 21496 26114 21548
rect 24636 21440 25176 21468
rect 24636 21428 24642 21440
rect 21358 21400 21364 21412
rect 20348 21372 21364 21400
rect 21358 21360 21364 21372
rect 21416 21360 21422 21412
rect 3421 21335 3479 21341
rect 3421 21301 3433 21335
rect 3467 21332 3479 21335
rect 3510 21332 3516 21344
rect 3467 21304 3516 21332
rect 3467 21301 3479 21304
rect 3421 21295 3479 21301
rect 3510 21292 3516 21304
rect 3568 21332 3574 21344
rect 3970 21332 3976 21344
rect 3568 21304 3976 21332
rect 3568 21292 3574 21304
rect 3970 21292 3976 21304
rect 4028 21292 4034 21344
rect 5626 21292 5632 21344
rect 5684 21292 5690 21344
rect 5718 21292 5724 21344
rect 5776 21292 5782 21344
rect 6178 21292 6184 21344
rect 6236 21292 6242 21344
rect 6638 21292 6644 21344
rect 6696 21332 6702 21344
rect 15562 21332 15568 21344
rect 6696 21304 15568 21332
rect 6696 21292 6702 21304
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 15654 21292 15660 21344
rect 15712 21292 15718 21344
rect 20162 21292 20168 21344
rect 20220 21332 20226 21344
rect 20806 21332 20812 21344
rect 20220 21304 20812 21332
rect 20220 21292 20226 21304
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 21910 21292 21916 21344
rect 21968 21292 21974 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24397 21335 24455 21341
rect 24397 21332 24409 21335
rect 24268 21304 24409 21332
rect 24268 21292 24274 21304
rect 24397 21301 24409 21304
rect 24443 21301 24455 21335
rect 24397 21295 24455 21301
rect 24765 21335 24823 21341
rect 24765 21301 24777 21335
rect 24811 21332 24823 21335
rect 24946 21332 24952 21344
rect 24811 21304 24952 21332
rect 24811 21301 24823 21304
rect 24765 21295 24823 21301
rect 24946 21292 24952 21304
rect 25004 21292 25010 21344
rect 25041 21335 25099 21341
rect 25041 21301 25053 21335
rect 25087 21332 25099 21335
rect 25498 21332 25504 21344
rect 25087 21304 25504 21332
rect 25087 21301 25099 21304
rect 25041 21295 25099 21301
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 25682 21292 25688 21344
rect 25740 21292 25746 21344
rect 1104 21242 26864 21264
rect 1104 21190 2918 21242
rect 2970 21190 2982 21242
rect 3034 21190 3046 21242
rect 3098 21190 3110 21242
rect 3162 21190 3174 21242
rect 3226 21190 3238 21242
rect 3290 21190 6918 21242
rect 6970 21190 6982 21242
rect 7034 21190 7046 21242
rect 7098 21190 7110 21242
rect 7162 21190 7174 21242
rect 7226 21190 7238 21242
rect 7290 21190 10918 21242
rect 10970 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 11238 21242
rect 11290 21190 14918 21242
rect 14970 21190 14982 21242
rect 15034 21190 15046 21242
rect 15098 21190 15110 21242
rect 15162 21190 15174 21242
rect 15226 21190 15238 21242
rect 15290 21190 18918 21242
rect 18970 21190 18982 21242
rect 19034 21190 19046 21242
rect 19098 21190 19110 21242
rect 19162 21190 19174 21242
rect 19226 21190 19238 21242
rect 19290 21190 22918 21242
rect 22970 21190 22982 21242
rect 23034 21190 23046 21242
rect 23098 21190 23110 21242
rect 23162 21190 23174 21242
rect 23226 21190 23238 21242
rect 23290 21190 26864 21242
rect 1104 21168 26864 21190
rect 2682 21088 2688 21140
rect 2740 21128 2746 21140
rect 3789 21131 3847 21137
rect 3789 21128 3801 21131
rect 2740 21100 3801 21128
rect 2740 21088 2746 21100
rect 3789 21097 3801 21100
rect 3835 21097 3847 21131
rect 3789 21091 3847 21097
rect 4430 21088 4436 21140
rect 4488 21128 4494 21140
rect 8202 21128 8208 21140
rect 4488 21100 8208 21128
rect 4488 21088 4494 21100
rect 8202 21088 8208 21100
rect 8260 21088 8266 21140
rect 10045 21131 10103 21137
rect 10045 21097 10057 21131
rect 10091 21128 10103 21131
rect 10226 21128 10232 21140
rect 10091 21100 10232 21128
rect 10091 21097 10103 21100
rect 10045 21091 10103 21097
rect 10226 21088 10232 21100
rect 10284 21088 10290 21140
rect 14458 21088 14464 21140
rect 14516 21128 14522 21140
rect 14553 21131 14611 21137
rect 14553 21128 14565 21131
rect 14516 21100 14565 21128
rect 14516 21088 14522 21100
rect 14553 21097 14565 21100
rect 14599 21097 14611 21131
rect 19610 21128 19616 21140
rect 14553 21091 14611 21097
rect 16868 21100 19616 21128
rect 1946 20952 1952 21004
rect 2004 20952 2010 21004
rect 4448 21001 4476 21088
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 5261 20995 5319 21001
rect 5261 20961 5273 20995
rect 5307 20992 5319 20995
rect 6454 20992 6460 21004
rect 5307 20964 6460 20992
rect 5307 20961 5319 20964
rect 5261 20955 5319 20961
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 16868 20992 16896 21100
rect 19610 21088 19616 21100
rect 19668 21088 19674 21140
rect 24762 21088 24768 21140
rect 24820 21088 24826 21140
rect 18506 21020 18512 21072
rect 18564 21060 18570 21072
rect 22094 21060 22100 21072
rect 18564 21032 19288 21060
rect 18564 21020 18570 21032
rect 12406 20964 16896 20992
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 4157 20927 4215 20933
rect 4157 20924 4169 20927
rect 4028 20896 4169 20924
rect 4028 20884 4034 20896
rect 4157 20893 4169 20896
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 5718 20884 5724 20936
rect 5776 20924 5782 20936
rect 9493 20927 9551 20933
rect 9493 20924 9505 20927
rect 5776 20896 9505 20924
rect 5776 20884 5782 20896
rect 9493 20893 9505 20896
rect 9539 20893 9551 20927
rect 9493 20887 9551 20893
rect 9582 20884 9588 20936
rect 9640 20884 9646 20936
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 9861 20927 9919 20933
rect 9861 20893 9873 20927
rect 9907 20924 9919 20927
rect 12406 20924 12434 20964
rect 9907 20896 12434 20924
rect 14737 20927 14795 20933
rect 9907 20893 9919 20896
rect 9861 20887 9919 20893
rect 14737 20893 14749 20927
rect 14783 20924 14795 20927
rect 15654 20924 15660 20936
rect 14783 20896 15660 20924
rect 14783 20893 14795 20896
rect 14737 20887 14795 20893
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 16942 20884 16948 20936
rect 17000 20884 17006 20936
rect 17126 20884 17132 20936
rect 17184 20884 17190 20936
rect 17586 20884 17592 20936
rect 17644 20884 17650 20936
rect 18322 20884 18328 20936
rect 18380 20884 18386 20936
rect 18598 20884 18604 20936
rect 18656 20884 18662 20936
rect 19260 20924 19288 21032
rect 22020 21032 22100 21060
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 22020 21001 22048 21032
rect 22094 21020 22100 21032
rect 22152 21020 22158 21072
rect 22005 20995 22063 21001
rect 19484 20964 19840 20992
rect 19484 20952 19490 20964
rect 19812 20933 19840 20964
rect 22005 20961 22017 20995
rect 22051 20992 22063 20995
rect 26513 20995 26571 21001
rect 26513 20992 26525 20995
rect 22051 20964 26525 20992
rect 22051 20961 22063 20964
rect 22005 20955 22063 20961
rect 26513 20961 26525 20964
rect 26559 20961 26571 20995
rect 26513 20955 26571 20961
rect 19337 20927 19395 20933
rect 19337 20924 19349 20927
rect 19260 20896 19349 20924
rect 19337 20893 19349 20896
rect 19383 20893 19395 20927
rect 19337 20887 19395 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 2216 20859 2274 20865
rect 2216 20825 2228 20859
rect 2262 20856 2274 20859
rect 2406 20856 2412 20868
rect 2262 20828 2412 20856
rect 2262 20825 2274 20828
rect 2216 20819 2274 20825
rect 2406 20816 2412 20828
rect 2464 20816 2470 20868
rect 5534 20816 5540 20868
rect 5592 20856 5598 20868
rect 6730 20865 6736 20868
rect 5997 20859 6055 20865
rect 5997 20856 6009 20859
rect 5592 20828 6009 20856
rect 5592 20816 5598 20828
rect 5997 20825 6009 20828
rect 6043 20825 6055 20859
rect 5997 20819 6055 20825
rect 6724 20819 6736 20865
rect 6730 20816 6736 20819
rect 6788 20816 6794 20868
rect 17144 20856 17172 20884
rect 18138 20856 18144 20868
rect 17144 20828 18144 20856
rect 18138 20816 18144 20828
rect 18196 20816 18202 20868
rect 18782 20816 18788 20868
rect 18840 20856 18846 20868
rect 19429 20859 19487 20865
rect 19429 20856 19441 20859
rect 18840 20828 19441 20856
rect 18840 20816 18846 20828
rect 19429 20825 19441 20828
rect 19475 20825 19487 20859
rect 19429 20819 19487 20825
rect 19518 20816 19524 20868
rect 19576 20856 19582 20868
rect 19904 20856 19932 20887
rect 20254 20884 20260 20936
rect 20312 20884 20318 20936
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20893 22155 20927
rect 22097 20887 22155 20893
rect 19576 20828 19932 20856
rect 19981 20859 20039 20865
rect 19576 20816 19582 20828
rect 19981 20825 19993 20859
rect 20027 20825 20039 20859
rect 19981 20819 20039 20825
rect 3326 20748 3332 20800
rect 3384 20748 3390 20800
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 4249 20791 4307 20797
rect 4249 20788 4261 20791
rect 4212 20760 4261 20788
rect 4212 20748 4218 20760
rect 4249 20757 4261 20760
rect 4295 20788 4307 20791
rect 5810 20788 5816 20800
rect 4295 20760 5816 20788
rect 4295 20757 4307 20760
rect 4249 20751 4307 20757
rect 5810 20748 5816 20760
rect 5868 20748 5874 20800
rect 7374 20748 7380 20800
rect 7432 20788 7438 20800
rect 7837 20791 7895 20797
rect 7837 20788 7849 20791
rect 7432 20760 7849 20788
rect 7432 20748 7438 20760
rect 7837 20757 7849 20760
rect 7883 20757 7895 20791
rect 7837 20751 7895 20757
rect 8754 20748 8760 20800
rect 8812 20788 8818 20800
rect 15562 20788 15568 20800
rect 8812 20760 15568 20788
rect 8812 20748 8818 20760
rect 15562 20748 15568 20760
rect 15620 20788 15626 20800
rect 16761 20791 16819 20797
rect 16761 20788 16773 20791
rect 15620 20760 16773 20788
rect 15620 20748 15626 20760
rect 16761 20757 16773 20760
rect 16807 20757 16819 20791
rect 18156 20788 18184 20816
rect 18690 20788 18696 20800
rect 18156 20760 18696 20788
rect 16761 20751 16819 20757
rect 18690 20748 18696 20760
rect 18748 20788 18754 20800
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 18748 20760 18889 20788
rect 18748 20748 18754 20760
rect 18877 20757 18889 20760
rect 18923 20788 18935 20791
rect 19996 20788 20024 20819
rect 18923 20760 20024 20788
rect 18923 20757 18935 20760
rect 18877 20751 18935 20757
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 22112 20788 22140 20887
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 23569 20927 23627 20933
rect 23569 20924 23581 20927
rect 23532 20896 23581 20924
rect 23532 20884 23538 20896
rect 23569 20893 23581 20896
rect 23615 20893 23627 20927
rect 23569 20887 23627 20893
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20924 23995 20927
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 23983 20896 24593 20924
rect 23983 20893 23995 20896
rect 23937 20887 23995 20893
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24673 20927 24731 20933
rect 24673 20893 24685 20927
rect 24719 20924 24731 20927
rect 24762 20924 24768 20936
rect 24719 20896 24768 20924
rect 24719 20893 24731 20896
rect 24673 20887 24731 20893
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 23753 20859 23811 20865
rect 23753 20825 23765 20859
rect 23799 20825 23811 20859
rect 23753 20819 23811 20825
rect 23845 20859 23903 20865
rect 23845 20825 23857 20859
rect 23891 20856 23903 20859
rect 24210 20856 24216 20868
rect 23891 20828 24216 20856
rect 23891 20825 23903 20828
rect 23845 20819 23903 20825
rect 20496 20760 22140 20788
rect 20496 20748 20502 20760
rect 22186 20748 22192 20800
rect 22244 20748 22250 20800
rect 23566 20748 23572 20800
rect 23624 20788 23630 20800
rect 23768 20788 23796 20819
rect 24210 20816 24216 20828
rect 24268 20816 24274 20868
rect 25682 20816 25688 20868
rect 25740 20816 25746 20868
rect 26142 20816 26148 20868
rect 26200 20856 26206 20868
rect 26237 20859 26295 20865
rect 26237 20856 26249 20859
rect 26200 20828 26249 20856
rect 26200 20816 26206 20828
rect 26237 20825 26249 20828
rect 26283 20825 26295 20859
rect 26237 20819 26295 20825
rect 23624 20760 23796 20788
rect 23624 20748 23630 20760
rect 24118 20748 24124 20800
rect 24176 20748 24182 20800
rect 1104 20698 26864 20720
rect 1104 20646 3658 20698
rect 3710 20646 3722 20698
rect 3774 20646 3786 20698
rect 3838 20646 3850 20698
rect 3902 20646 3914 20698
rect 3966 20646 3978 20698
rect 4030 20646 7658 20698
rect 7710 20646 7722 20698
rect 7774 20646 7786 20698
rect 7838 20646 7850 20698
rect 7902 20646 7914 20698
rect 7966 20646 7978 20698
rect 8030 20646 11658 20698
rect 11710 20646 11722 20698
rect 11774 20646 11786 20698
rect 11838 20646 11850 20698
rect 11902 20646 11914 20698
rect 11966 20646 11978 20698
rect 12030 20646 15658 20698
rect 15710 20646 15722 20698
rect 15774 20646 15786 20698
rect 15838 20646 15850 20698
rect 15902 20646 15914 20698
rect 15966 20646 15978 20698
rect 16030 20646 19658 20698
rect 19710 20646 19722 20698
rect 19774 20646 19786 20698
rect 19838 20646 19850 20698
rect 19902 20646 19914 20698
rect 19966 20646 19978 20698
rect 20030 20646 23658 20698
rect 23710 20646 23722 20698
rect 23774 20646 23786 20698
rect 23838 20646 23850 20698
rect 23902 20646 23914 20698
rect 23966 20646 23978 20698
rect 24030 20646 26864 20698
rect 1104 20624 26864 20646
rect 2406 20544 2412 20596
rect 2464 20544 2470 20596
rect 2869 20587 2927 20593
rect 2869 20584 2881 20587
rect 2746 20556 2881 20584
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20448 2651 20451
rect 2746 20448 2774 20556
rect 2869 20553 2881 20556
rect 2915 20553 2927 20587
rect 2869 20547 2927 20553
rect 3237 20587 3295 20593
rect 3237 20553 3249 20587
rect 3283 20584 3295 20587
rect 3326 20584 3332 20596
rect 3283 20556 3332 20584
rect 3283 20553 3295 20556
rect 3237 20547 3295 20553
rect 3326 20544 3332 20556
rect 3384 20544 3390 20596
rect 4890 20544 4896 20596
rect 4948 20544 4954 20596
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 5626 20584 5632 20596
rect 5307 20556 5632 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 6730 20544 6736 20596
rect 6788 20544 6794 20596
rect 7009 20587 7067 20593
rect 7009 20553 7021 20587
rect 7055 20553 7067 20587
rect 7009 20547 7067 20553
rect 2639 20420 2774 20448
rect 3344 20448 3372 20544
rect 3510 20476 3516 20528
rect 3568 20516 3574 20528
rect 4065 20519 4123 20525
rect 4065 20516 4077 20519
rect 3568 20488 4077 20516
rect 3568 20476 3574 20488
rect 4065 20485 4077 20488
rect 4111 20485 4123 20519
rect 4065 20479 4123 20485
rect 5353 20519 5411 20525
rect 5353 20485 5365 20519
rect 5399 20516 5411 20519
rect 5810 20516 5816 20528
rect 5399 20488 5816 20516
rect 5399 20485 5411 20488
rect 5353 20479 5411 20485
rect 5810 20476 5816 20488
rect 5868 20476 5874 20528
rect 3789 20451 3847 20457
rect 3789 20448 3801 20451
rect 3344 20420 3801 20448
rect 2639 20417 2651 20420
rect 2593 20411 2651 20417
rect 3789 20417 3801 20420
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 3970 20408 3976 20460
rect 4028 20408 4034 20460
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20448 4215 20451
rect 4246 20448 4252 20460
rect 4203 20420 4252 20448
rect 4203 20417 4215 20420
rect 4157 20411 4215 20417
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 5258 20408 5264 20460
rect 5316 20448 5322 20460
rect 6917 20451 6975 20457
rect 5316 20420 5488 20448
rect 5316 20408 5322 20420
rect 3329 20383 3387 20389
rect 3329 20349 3341 20383
rect 3375 20349 3387 20383
rect 3329 20343 3387 20349
rect 3344 20312 3372 20343
rect 3510 20340 3516 20392
rect 3568 20340 3574 20392
rect 5460 20389 5488 20420
rect 6917 20417 6929 20451
rect 6963 20448 6975 20451
rect 7024 20448 7052 20547
rect 7374 20544 7380 20596
rect 7432 20544 7438 20596
rect 7650 20544 7656 20596
rect 7708 20584 7714 20596
rect 12802 20584 12808 20596
rect 7708 20556 12808 20584
rect 7708 20544 7714 20556
rect 12802 20544 12808 20556
rect 12860 20584 12866 20596
rect 15378 20584 15384 20596
rect 12860 20556 15384 20584
rect 12860 20544 12866 20556
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 18598 20584 18604 20596
rect 17420 20556 18604 20584
rect 7469 20519 7527 20525
rect 7469 20485 7481 20519
rect 7515 20516 7527 20519
rect 8202 20516 8208 20528
rect 7515 20488 8208 20516
rect 7515 20485 7527 20488
rect 7469 20479 7527 20485
rect 8202 20476 8208 20488
rect 8260 20516 8266 20528
rect 9953 20519 10011 20525
rect 9953 20516 9965 20519
rect 8260 20488 9965 20516
rect 8260 20476 8266 20488
rect 9953 20485 9965 20488
rect 9999 20516 10011 20519
rect 12250 20516 12256 20528
rect 9999 20488 12256 20516
rect 9999 20485 10011 20488
rect 9953 20479 10011 20485
rect 12250 20476 12256 20488
rect 12308 20476 12314 20528
rect 14093 20519 14151 20525
rect 14093 20485 14105 20519
rect 14139 20516 14151 20519
rect 16482 20516 16488 20528
rect 14139 20488 16488 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 9861 20451 9919 20457
rect 6963 20420 7052 20448
rect 7116 20420 7604 20448
rect 6963 20417 6975 20420
rect 6917 20411 6975 20417
rect 5445 20383 5503 20389
rect 5445 20349 5457 20383
rect 5491 20380 5503 20383
rect 7116 20380 7144 20420
rect 7576 20389 7604 20420
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10318 20448 10324 20460
rect 9907 20420 10324 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 13262 20408 13268 20460
rect 13320 20408 13326 20460
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 13722 20408 13728 20460
rect 13780 20448 13786 20460
rect 13998 20457 14004 20460
rect 13817 20451 13875 20457
rect 13817 20448 13829 20451
rect 13780 20420 13829 20448
rect 13780 20408 13786 20420
rect 13817 20417 13829 20420
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 13965 20451 14004 20457
rect 13965 20417 13977 20451
rect 13965 20411 14004 20417
rect 13998 20408 14004 20411
rect 14056 20408 14062 20460
rect 5491 20352 7144 20380
rect 7561 20383 7619 20389
rect 5491 20349 5503 20352
rect 5445 20343 5503 20349
rect 7561 20349 7573 20383
rect 7607 20349 7619 20383
rect 7561 20343 7619 20349
rect 10042 20340 10048 20392
rect 10100 20380 10106 20392
rect 10137 20383 10195 20389
rect 10137 20380 10149 20383
rect 10100 20352 10149 20380
rect 10100 20340 10106 20352
rect 10137 20349 10149 20352
rect 10183 20380 10195 20383
rect 13446 20380 13452 20392
rect 10183 20352 13452 20380
rect 10183 20349 10195 20352
rect 10137 20343 10195 20349
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 4154 20312 4160 20324
rect 3344 20284 4160 20312
rect 4154 20272 4160 20284
rect 4212 20272 4218 20324
rect 4341 20315 4399 20321
rect 4341 20281 4353 20315
rect 4387 20312 4399 20315
rect 6362 20312 6368 20324
rect 4387 20284 6368 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 6362 20272 6368 20284
rect 6420 20272 6426 20324
rect 14108 20312 14136 20479
rect 16482 20476 16488 20488
rect 16540 20476 16546 20528
rect 17420 20525 17448 20556
rect 18598 20544 18604 20556
rect 18656 20584 18662 20596
rect 18656 20556 18828 20584
rect 18656 20544 18662 20556
rect 17405 20519 17463 20525
rect 17405 20485 17417 20519
rect 17451 20485 17463 20519
rect 17405 20479 17463 20485
rect 17957 20519 18015 20525
rect 17957 20485 17969 20519
rect 18003 20516 18015 20519
rect 18322 20516 18328 20528
rect 18003 20488 18328 20516
rect 18003 20485 18015 20488
rect 17957 20479 18015 20485
rect 18322 20476 18328 20488
rect 18380 20516 18386 20528
rect 18800 20525 18828 20556
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20312 20556 21097 20584
rect 20312 20544 20318 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 21453 20587 21511 20593
rect 21453 20553 21465 20587
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 24029 20587 24087 20593
rect 24029 20553 24041 20587
rect 24075 20553 24087 20587
rect 24029 20547 24087 20553
rect 18785 20519 18843 20525
rect 18380 20488 18736 20516
rect 18380 20476 18386 20488
rect 18708 20460 18736 20488
rect 18785 20485 18797 20519
rect 18831 20516 18843 20519
rect 19518 20516 19524 20528
rect 18831 20488 19524 20516
rect 18831 20485 18843 20488
rect 18785 20479 18843 20485
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 19610 20476 19616 20528
rect 19668 20516 19674 20528
rect 19668 20488 20300 20516
rect 19668 20476 19674 20488
rect 14366 20457 14372 20460
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 14323 20451 14372 20457
rect 14323 20417 14335 20451
rect 14369 20417 14372 20451
rect 14323 20411 14372 20417
rect 14200 20380 14228 20411
rect 14366 20408 14372 20411
rect 14424 20448 14430 20460
rect 17497 20451 17555 20457
rect 14424 20420 16528 20448
rect 14424 20408 14430 20420
rect 14200 20352 14320 20380
rect 14292 20324 14320 20352
rect 6472 20284 14136 20312
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 6472 20244 6500 20284
rect 14274 20272 14280 20324
rect 14332 20272 14338 20324
rect 4028 20216 6500 20244
rect 4028 20204 4034 20216
rect 8570 20204 8576 20256
rect 8628 20244 8634 20256
rect 9493 20247 9551 20253
rect 9493 20244 9505 20247
rect 8628 20216 9505 20244
rect 8628 20204 8634 20216
rect 9493 20213 9505 20216
rect 9539 20213 9551 20247
rect 9493 20207 9551 20213
rect 13078 20204 13084 20256
rect 13136 20204 13142 20256
rect 13354 20204 13360 20256
rect 13412 20204 13418 20256
rect 13906 20204 13912 20256
rect 13964 20244 13970 20256
rect 14461 20247 14519 20253
rect 14461 20244 14473 20247
rect 13964 20216 14473 20244
rect 13964 20204 13970 20216
rect 14461 20213 14473 20216
rect 14507 20213 14519 20247
rect 16500 20244 16528 20420
rect 17497 20417 17509 20451
rect 17543 20448 17555 20451
rect 18506 20448 18512 20460
rect 17543 20420 18512 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 18506 20408 18512 20420
rect 18564 20408 18570 20460
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 19334 20448 19340 20460
rect 18748 20420 19340 20448
rect 18748 20408 18754 20420
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 19429 20451 19487 20457
rect 19429 20417 19441 20451
rect 19475 20448 19487 20451
rect 19475 20420 19840 20448
rect 19475 20417 19487 20420
rect 19429 20411 19487 20417
rect 19812 20392 19840 20420
rect 19886 20408 19892 20460
rect 19944 20408 19950 20460
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20162 20448 20168 20460
rect 20027 20420 20168 20448
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20272 20457 20300 20488
rect 20438 20476 20444 20528
rect 20496 20476 20502 20528
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20714 20448 20720 20460
rect 20303 20420 20720 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 21468 20448 21496 20547
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21468 20420 21833 20448
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 22646 20408 22652 20460
rect 22704 20408 22710 20460
rect 23569 20451 23627 20457
rect 23569 20417 23581 20451
rect 23615 20417 23627 20451
rect 24044 20448 24072 20547
rect 24394 20544 24400 20596
rect 24452 20584 24458 20596
rect 24765 20587 24823 20593
rect 24765 20584 24777 20587
rect 24452 20556 24777 20584
rect 24452 20544 24458 20556
rect 24765 20553 24777 20556
rect 24811 20553 24823 20587
rect 24765 20547 24823 20553
rect 24946 20544 24952 20596
rect 25004 20584 25010 20596
rect 25133 20587 25191 20593
rect 25133 20584 25145 20587
rect 25004 20556 25145 20584
rect 25004 20544 25010 20556
rect 25133 20553 25145 20556
rect 25179 20553 25191 20587
rect 25133 20547 25191 20553
rect 24118 20476 24124 20528
rect 24176 20476 24182 20528
rect 25041 20451 25099 20457
rect 25041 20448 25053 20451
rect 24044 20420 25053 20448
rect 23569 20411 23627 20417
rect 25041 20417 25053 20420
rect 25087 20417 25099 20451
rect 25041 20411 25099 20417
rect 16942 20340 16948 20392
rect 17000 20340 17006 20392
rect 17862 20340 17868 20392
rect 17920 20340 17926 20392
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 18233 20383 18291 20389
rect 18233 20380 18245 20383
rect 18196 20352 18245 20380
rect 18196 20340 18202 20352
rect 18233 20349 18245 20352
rect 18279 20349 18291 20383
rect 18233 20343 18291 20349
rect 18322 20340 18328 20392
rect 18380 20340 18386 20392
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 19245 20383 19303 20389
rect 19245 20380 19257 20383
rect 18472 20352 19257 20380
rect 18472 20340 18478 20352
rect 19245 20349 19257 20352
rect 19291 20349 19303 20383
rect 19245 20343 19303 20349
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19702 20380 19708 20392
rect 19567 20352 19708 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19702 20340 19708 20352
rect 19760 20340 19766 20392
rect 19794 20340 19800 20392
rect 19852 20380 19858 20392
rect 20346 20380 20352 20392
rect 19852 20352 20352 20380
rect 19852 20340 19858 20352
rect 20346 20340 20352 20352
rect 20404 20340 20410 20392
rect 20898 20340 20904 20392
rect 20956 20340 20962 20392
rect 20993 20383 21051 20389
rect 20993 20349 21005 20383
rect 21039 20380 21051 20383
rect 22186 20380 22192 20392
rect 21039 20352 22192 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 22186 20340 22192 20352
rect 22244 20340 22250 20392
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20380 22523 20383
rect 22554 20380 22560 20392
rect 22511 20352 22560 20380
rect 22511 20349 22523 20352
rect 22465 20343 22523 20349
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 23584 20380 23612 20411
rect 25498 20408 25504 20460
rect 25556 20408 25562 20460
rect 25774 20408 25780 20460
rect 25832 20448 25838 20460
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 25832 20420 26065 20448
rect 25832 20408 25838 20420
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 24118 20380 24124 20392
rect 23584 20352 24124 20380
rect 24118 20340 24124 20352
rect 24176 20340 24182 20392
rect 24489 20383 24547 20389
rect 24489 20349 24501 20383
rect 24535 20380 24547 20383
rect 24670 20380 24676 20392
rect 24535 20352 24676 20380
rect 24535 20349 24547 20352
rect 24489 20343 24547 20349
rect 24670 20340 24676 20352
rect 24728 20340 24734 20392
rect 25225 20383 25283 20389
rect 25225 20349 25237 20383
rect 25271 20349 25283 20383
rect 25225 20343 25283 20349
rect 25409 20383 25467 20389
rect 25409 20349 25421 20383
rect 25455 20380 25467 20383
rect 26418 20380 26424 20392
rect 25455 20352 26424 20380
rect 25455 20349 25467 20352
rect 25409 20343 25467 20349
rect 16960 20312 16988 20340
rect 18432 20312 18460 20340
rect 16960 20284 18460 20312
rect 24286 20315 24344 20321
rect 24286 20281 24298 20315
rect 24332 20312 24344 20315
rect 24949 20315 25007 20321
rect 24949 20312 24961 20315
rect 24332 20284 24961 20312
rect 24332 20281 24344 20284
rect 24286 20275 24344 20281
rect 24949 20281 24961 20284
rect 24995 20281 25007 20315
rect 25240 20312 25268 20343
rect 26418 20340 26424 20352
rect 26476 20340 26482 20392
rect 25593 20315 25651 20321
rect 25593 20312 25605 20315
rect 25240 20284 25605 20312
rect 24949 20275 25007 20281
rect 25593 20281 25605 20284
rect 25639 20281 25651 20315
rect 25593 20275 25651 20281
rect 18782 20244 18788 20256
rect 16500 20216 18788 20244
rect 14461 20207 14519 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 20530 20244 20536 20256
rect 19576 20216 20536 20244
rect 19576 20204 19582 20216
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 22002 20204 22008 20256
rect 22060 20204 22066 20256
rect 23474 20204 23480 20256
rect 23532 20244 23538 20256
rect 23658 20244 23664 20256
rect 23532 20216 23664 20244
rect 23532 20204 23538 20216
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 24394 20204 24400 20256
rect 24452 20204 24458 20256
rect 25222 20204 25228 20256
rect 25280 20244 25286 20256
rect 25777 20247 25835 20253
rect 25777 20244 25789 20247
rect 25280 20216 25789 20244
rect 25280 20204 25286 20216
rect 25777 20213 25789 20216
rect 25823 20213 25835 20247
rect 25777 20207 25835 20213
rect 1104 20154 26864 20176
rect 1104 20102 2918 20154
rect 2970 20102 2982 20154
rect 3034 20102 3046 20154
rect 3098 20102 3110 20154
rect 3162 20102 3174 20154
rect 3226 20102 3238 20154
rect 3290 20102 6918 20154
rect 6970 20102 6982 20154
rect 7034 20102 7046 20154
rect 7098 20102 7110 20154
rect 7162 20102 7174 20154
rect 7226 20102 7238 20154
rect 7290 20102 10918 20154
rect 10970 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 11238 20154
rect 11290 20102 14918 20154
rect 14970 20102 14982 20154
rect 15034 20102 15046 20154
rect 15098 20102 15110 20154
rect 15162 20102 15174 20154
rect 15226 20102 15238 20154
rect 15290 20102 18918 20154
rect 18970 20102 18982 20154
rect 19034 20102 19046 20154
rect 19098 20102 19110 20154
rect 19162 20102 19174 20154
rect 19226 20102 19238 20154
rect 19290 20102 22918 20154
rect 22970 20102 22982 20154
rect 23034 20102 23046 20154
rect 23098 20102 23110 20154
rect 23162 20102 23174 20154
rect 23226 20102 23238 20154
rect 23290 20102 26864 20154
rect 1104 20080 26864 20102
rect 5166 20040 5172 20052
rect 4632 20012 5172 20040
rect 3329 19975 3387 19981
rect 3329 19941 3341 19975
rect 3375 19941 3387 19975
rect 3329 19935 3387 19941
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19836 2007 19839
rect 2498 19836 2504 19848
rect 1995 19808 2504 19836
rect 1995 19805 2007 19808
rect 1949 19799 2007 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 3142 19796 3148 19848
rect 3200 19836 3206 19848
rect 3344 19836 3372 19935
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 3200 19808 3801 19836
rect 3200 19796 3206 19808
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 3970 19796 3976 19848
rect 4028 19796 4034 19848
rect 4062 19796 4068 19848
rect 4120 19796 4126 19848
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4632 19836 4660 20012
rect 5166 20000 5172 20012
rect 5224 20040 5230 20052
rect 7006 20040 7012 20052
rect 5224 20012 7012 20040
rect 5224 20000 5230 20012
rect 7006 20000 7012 20012
rect 7064 20040 7070 20052
rect 7650 20040 7656 20052
rect 7064 20012 7656 20040
rect 7064 20000 7070 20012
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 13262 20000 13268 20052
rect 13320 20040 13326 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13320 20012 14105 20040
rect 13320 20000 13326 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 19245 20043 19303 20049
rect 19245 20040 19257 20043
rect 14093 20003 14151 20009
rect 14200 20012 19257 20040
rect 13722 19932 13728 19984
rect 13780 19972 13786 19984
rect 14200 19972 14228 20012
rect 19245 20009 19257 20012
rect 19291 20009 19303 20043
rect 19245 20003 19303 20009
rect 20254 20000 20260 20052
rect 20312 20040 20318 20052
rect 20312 20012 22600 20040
rect 20312 20000 20318 20012
rect 13780 19944 14228 19972
rect 17926 19944 18276 19972
rect 13780 19932 13786 19944
rect 8662 19864 8668 19916
rect 8720 19904 8726 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 8720 19876 8953 19904
rect 8720 19864 8726 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 8941 19867 8999 19873
rect 4203 19808 4660 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 6638 19836 6644 19848
rect 4764 19808 6644 19836
rect 4764 19796 4770 19808
rect 6638 19796 6644 19808
rect 6696 19836 6702 19848
rect 6733 19839 6791 19845
rect 6733 19836 6745 19839
rect 6696 19808 6745 19836
rect 6696 19796 6702 19808
rect 6733 19805 6745 19808
rect 6779 19805 6791 19839
rect 6733 19799 6791 19805
rect 8570 19796 8576 19848
rect 8628 19796 8634 19848
rect 8956 19836 8984 19867
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 14645 19907 14703 19913
rect 14645 19904 14657 19907
rect 14240 19876 14657 19904
rect 14240 19864 14246 19876
rect 14645 19873 14657 19876
rect 14691 19873 14703 19907
rect 16942 19904 16948 19916
rect 14645 19867 14703 19873
rect 16316 19876 16948 19904
rect 10597 19839 10655 19845
rect 10597 19836 10609 19839
rect 8956 19808 10609 19836
rect 10597 19805 10609 19808
rect 10643 19836 10655 19839
rect 10962 19836 10968 19848
rect 10643 19808 10968 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 10962 19796 10968 19808
rect 11020 19836 11026 19848
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 11020 19808 11069 19836
rect 11020 19796 11026 19808
rect 11057 19805 11069 19808
rect 11103 19836 11115 19839
rect 12526 19836 12532 19848
rect 11103 19808 12532 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12796 19839 12854 19845
rect 12796 19805 12808 19839
rect 12842 19836 12854 19839
rect 13354 19836 13360 19848
rect 12842 19808 13360 19836
rect 12842 19805 12854 19808
rect 12796 19799 12854 19805
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 16316 19845 16344 19876
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17926 19904 17954 19944
rect 18049 19907 18107 19913
rect 18049 19904 18061 19907
rect 17052 19876 18061 19904
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 14056 19808 14473 19836
rect 14056 19796 14062 19808
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 16758 19796 16764 19848
rect 16816 19836 16822 19848
rect 17052 19845 17080 19876
rect 18049 19873 18061 19876
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 18138 19864 18144 19916
rect 18196 19864 18202 19916
rect 18248 19904 18276 19944
rect 18966 19904 18972 19916
rect 18248 19876 18972 19904
rect 18966 19864 18972 19876
rect 19024 19904 19030 19916
rect 19610 19904 19616 19916
rect 19024 19876 19616 19904
rect 19024 19864 19030 19876
rect 19610 19864 19616 19876
rect 19668 19864 19674 19916
rect 19702 19864 19708 19916
rect 19760 19904 19766 19916
rect 20346 19904 20352 19916
rect 19760 19876 20352 19904
rect 19760 19864 19766 19876
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 22002 19864 22008 19916
rect 22060 19864 22066 19916
rect 22462 19864 22468 19916
rect 22520 19864 22526 19916
rect 17037 19839 17095 19845
rect 17037 19836 17049 19839
rect 16816 19808 17049 19836
rect 16816 19796 16822 19808
rect 17037 19805 17049 19808
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19836 17463 19839
rect 17586 19836 17592 19848
rect 17451 19808 17592 19836
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 18156 19836 18184 19864
rect 17828 19808 18184 19836
rect 17828 19796 17834 19808
rect 18506 19796 18512 19848
rect 18564 19796 18570 19848
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19805 19119 19839
rect 19061 19799 19119 19805
rect 2216 19771 2274 19777
rect 2216 19737 2228 19771
rect 2262 19768 2274 19771
rect 2406 19768 2412 19780
rect 2262 19740 2412 19768
rect 2262 19737 2274 19740
rect 2216 19731 2274 19737
rect 2406 19728 2412 19740
rect 2464 19728 2470 19780
rect 6546 19728 6552 19780
rect 6604 19768 6610 19780
rect 6978 19771 7036 19777
rect 6978 19768 6990 19771
rect 6604 19740 6990 19768
rect 6604 19728 6610 19740
rect 6978 19737 6990 19740
rect 7024 19737 7036 19771
rect 9186 19771 9244 19777
rect 9186 19768 9198 19771
rect 6978 19731 7036 19737
rect 8772 19740 9198 19768
rect 4341 19703 4399 19709
rect 4341 19669 4353 19703
rect 4387 19700 4399 19703
rect 4798 19700 4804 19712
rect 4387 19672 4804 19700
rect 4387 19669 4399 19672
rect 4341 19663 4399 19669
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 6086 19660 6092 19712
rect 6144 19700 6150 19712
rect 6730 19700 6736 19712
rect 6144 19672 6736 19700
rect 6144 19660 6150 19672
rect 6730 19660 6736 19672
rect 6788 19700 6794 19712
rect 7190 19700 7196 19712
rect 6788 19672 7196 19700
rect 6788 19660 6794 19672
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 8110 19660 8116 19712
rect 8168 19660 8174 19712
rect 8772 19709 8800 19740
rect 9186 19737 9198 19740
rect 9232 19737 9244 19771
rect 9186 19731 9244 19737
rect 11324 19771 11382 19777
rect 11324 19737 11336 19771
rect 11370 19768 11382 19771
rect 11514 19768 11520 19780
rect 11370 19740 11520 19768
rect 11370 19737 11382 19740
rect 11324 19731 11382 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 13630 19768 13636 19780
rect 13372 19740 13636 19768
rect 13372 19712 13400 19740
rect 13630 19728 13636 19740
rect 13688 19768 13694 19780
rect 14553 19771 14611 19777
rect 14553 19768 14565 19771
rect 13688 19740 14565 19768
rect 13688 19728 13694 19740
rect 14553 19737 14565 19740
rect 14599 19768 14611 19771
rect 14642 19768 14648 19780
rect 14599 19740 14648 19768
rect 14599 19737 14611 19740
rect 14553 19731 14611 19737
rect 14642 19728 14648 19740
rect 14700 19728 14706 19780
rect 18141 19771 18199 19777
rect 18141 19737 18153 19771
rect 18187 19768 18199 19771
rect 18322 19768 18328 19780
rect 18187 19740 18328 19768
rect 18187 19737 18199 19740
rect 18141 19731 18199 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 18414 19728 18420 19780
rect 18472 19768 18478 19780
rect 18601 19771 18659 19777
rect 18601 19768 18613 19771
rect 18472 19740 18613 19768
rect 18472 19728 18478 19740
rect 18601 19737 18613 19740
rect 18647 19737 18659 19771
rect 18601 19731 18659 19737
rect 19076 19768 19104 19799
rect 19518 19796 19524 19848
rect 19576 19796 19582 19848
rect 19794 19796 19800 19848
rect 19852 19796 19858 19848
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 22572 19845 22600 20012
rect 23566 20000 23572 20052
rect 23624 20040 23630 20052
rect 24029 20043 24087 20049
rect 24029 20040 24041 20043
rect 23624 20012 24041 20040
rect 23624 20000 23630 20012
rect 24029 20009 24041 20012
rect 24075 20009 24087 20043
rect 24029 20003 24087 20009
rect 24670 20000 24676 20052
rect 24728 20000 24734 20052
rect 22925 19975 22983 19981
rect 22925 19941 22937 19975
rect 22971 19972 22983 19975
rect 24394 19972 24400 19984
rect 22971 19944 24400 19972
rect 22971 19941 22983 19944
rect 22925 19935 22983 19941
rect 24394 19932 24400 19944
rect 24452 19932 24458 19984
rect 25498 19932 25504 19984
rect 25556 19932 25562 19984
rect 25516 19904 25544 19932
rect 24964 19876 25544 19904
rect 22281 19839 22339 19845
rect 22281 19805 22293 19839
rect 22327 19805 22339 19839
rect 22281 19799 22339 19805
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 23937 19839 23995 19845
rect 23937 19805 23949 19839
rect 23983 19836 23995 19839
rect 24118 19836 24124 19848
rect 23983 19808 24124 19836
rect 23983 19805 23995 19808
rect 23937 19799 23995 19805
rect 19334 19768 19340 19780
rect 19076 19740 19340 19768
rect 8757 19703 8815 19709
rect 8757 19669 8769 19703
rect 8803 19669 8815 19703
rect 8757 19663 8815 19669
rect 10318 19660 10324 19712
rect 10376 19660 10382 19712
rect 12158 19660 12164 19712
rect 12216 19700 12222 19712
rect 12437 19703 12495 19709
rect 12437 19700 12449 19703
rect 12216 19672 12449 19700
rect 12216 19660 12222 19672
rect 12437 19669 12449 19672
rect 12483 19669 12495 19703
rect 12437 19663 12495 19669
rect 13354 19660 13360 19712
rect 13412 19660 13418 19712
rect 13909 19703 13967 19709
rect 13909 19669 13921 19703
rect 13955 19700 13967 19703
rect 14274 19700 14280 19712
rect 13955 19672 14280 19700
rect 13955 19669 13967 19672
rect 13909 19663 13967 19669
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 16482 19660 16488 19712
rect 16540 19700 16546 19712
rect 16669 19703 16727 19709
rect 16669 19700 16681 19703
rect 16540 19672 16681 19700
rect 16540 19660 16546 19672
rect 16669 19669 16681 19672
rect 16715 19669 16727 19703
rect 16669 19663 16727 19669
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 19076 19700 19104 19740
rect 19334 19728 19340 19740
rect 19392 19768 19398 19780
rect 20438 19768 20444 19780
rect 19392 19740 20444 19768
rect 19392 19728 19398 19740
rect 20438 19728 20444 19740
rect 20496 19728 20502 19780
rect 21910 19768 21916 19780
rect 21574 19740 21916 19768
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 22094 19728 22100 19780
rect 22152 19768 22158 19780
rect 22296 19768 22324 19799
rect 24118 19796 24124 19808
rect 24176 19796 24182 19848
rect 24964 19845 24992 19876
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19805 24915 19839
rect 24857 19799 24915 19805
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 22152 19740 22324 19768
rect 24872 19768 24900 19799
rect 25222 19796 25228 19848
rect 25280 19796 25286 19848
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 25774 19836 25780 19848
rect 25547 19808 25780 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 25774 19796 25780 19808
rect 25832 19796 25838 19848
rect 25041 19771 25099 19777
rect 24872 19740 24992 19768
rect 22152 19728 22158 19740
rect 17644 19672 19104 19700
rect 17644 19660 17650 19672
rect 20254 19660 20260 19712
rect 20312 19700 20318 19712
rect 20533 19703 20591 19709
rect 20533 19700 20545 19703
rect 20312 19672 20545 19700
rect 20312 19660 20318 19672
rect 20533 19669 20545 19672
rect 20579 19669 20591 19703
rect 24964 19700 24992 19740
rect 25041 19737 25053 19771
rect 25087 19768 25099 19771
rect 25409 19771 25467 19777
rect 25409 19768 25421 19771
rect 25087 19740 25421 19768
rect 25087 19737 25099 19740
rect 25041 19731 25099 19737
rect 25409 19737 25421 19740
rect 25455 19737 25467 19771
rect 25409 19731 25467 19737
rect 26418 19700 26424 19712
rect 24964 19672 26424 19700
rect 20533 19663 20591 19669
rect 26418 19660 26424 19672
rect 26476 19660 26482 19712
rect 1104 19610 26864 19632
rect 1104 19558 3658 19610
rect 3710 19558 3722 19610
rect 3774 19558 3786 19610
rect 3838 19558 3850 19610
rect 3902 19558 3914 19610
rect 3966 19558 3978 19610
rect 4030 19558 7658 19610
rect 7710 19558 7722 19610
rect 7774 19558 7786 19610
rect 7838 19558 7850 19610
rect 7902 19558 7914 19610
rect 7966 19558 7978 19610
rect 8030 19558 11658 19610
rect 11710 19558 11722 19610
rect 11774 19558 11786 19610
rect 11838 19558 11850 19610
rect 11902 19558 11914 19610
rect 11966 19558 11978 19610
rect 12030 19558 15658 19610
rect 15710 19558 15722 19610
rect 15774 19558 15786 19610
rect 15838 19558 15850 19610
rect 15902 19558 15914 19610
rect 15966 19558 15978 19610
rect 16030 19558 19658 19610
rect 19710 19558 19722 19610
rect 19774 19558 19786 19610
rect 19838 19558 19850 19610
rect 19902 19558 19914 19610
rect 19966 19558 19978 19610
rect 20030 19558 23658 19610
rect 23710 19558 23722 19610
rect 23774 19558 23786 19610
rect 23838 19558 23850 19610
rect 23902 19558 23914 19610
rect 23966 19558 23978 19610
rect 24030 19558 26864 19610
rect 1104 19536 26864 19558
rect 2406 19456 2412 19508
rect 2464 19456 2470 19508
rect 2777 19499 2835 19505
rect 2777 19465 2789 19499
rect 2823 19465 2835 19499
rect 2777 19459 2835 19465
rect 2593 19363 2651 19369
rect 2593 19329 2605 19363
rect 2639 19360 2651 19363
rect 2792 19360 2820 19459
rect 3142 19456 3148 19508
rect 3200 19456 3206 19508
rect 6546 19456 6552 19508
rect 6604 19456 6610 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 6932 19468 7849 19496
rect 4062 19388 4068 19440
rect 4120 19428 4126 19440
rect 4706 19428 4712 19440
rect 4120 19400 4712 19428
rect 4120 19388 4126 19400
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 6454 19388 6460 19440
rect 6512 19428 6518 19440
rect 6512 19400 6776 19428
rect 6512 19388 6518 19400
rect 2639 19332 2820 19360
rect 3237 19363 3295 19369
rect 2639 19329 2651 19332
rect 2593 19323 2651 19329
rect 3237 19329 3249 19363
rect 3283 19360 3295 19363
rect 3326 19360 3332 19372
rect 3283 19332 3332 19360
rect 3283 19329 3295 19332
rect 3237 19323 3295 19329
rect 3326 19320 3332 19332
rect 3384 19360 3390 19372
rect 4246 19360 4252 19372
rect 3384 19332 4252 19360
rect 3384 19320 3390 19332
rect 4246 19320 4252 19332
rect 4304 19320 4310 19372
rect 5442 19320 5448 19372
rect 5500 19320 5506 19372
rect 6748 19369 6776 19400
rect 6932 19369 6960 19468
rect 7837 19465 7849 19468
rect 7883 19496 7895 19499
rect 8110 19496 8116 19508
rect 7883 19468 8116 19496
rect 7883 19465 7895 19468
rect 7837 19459 7895 19465
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 9401 19499 9459 19505
rect 9401 19465 9413 19499
rect 9447 19496 9459 19499
rect 10318 19496 10324 19508
rect 9447 19468 10324 19496
rect 9447 19465 9459 19468
rect 9401 19459 9459 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 10428 19468 11284 19496
rect 7006 19388 7012 19440
rect 7064 19388 7070 19440
rect 7098 19388 7104 19440
rect 7156 19388 7162 19440
rect 7374 19388 7380 19440
rect 7432 19428 7438 19440
rect 7432 19400 8340 19428
rect 7432 19388 7438 19400
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19360 6423 19363
rect 6733 19363 6791 19369
rect 6411 19332 6684 19360
rect 6411 19329 6423 19332
rect 6365 19323 6423 19329
rect 3421 19295 3479 19301
rect 3421 19261 3433 19295
rect 3467 19292 3479 19295
rect 3510 19292 3516 19304
rect 3467 19264 3516 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 3510 19252 3516 19264
rect 3568 19292 3574 19304
rect 6656 19292 6684 19332
rect 6733 19329 6745 19363
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 6881 19363 6960 19369
rect 6881 19329 6893 19363
rect 6927 19332 6960 19363
rect 6927 19329 6939 19332
rect 6881 19323 6939 19329
rect 7190 19320 7196 19372
rect 7248 19369 7254 19372
rect 7248 19360 7256 19369
rect 7929 19363 7987 19369
rect 7248 19332 7293 19360
rect 7248 19323 7256 19332
rect 7929 19329 7941 19363
rect 7975 19360 7987 19363
rect 8202 19360 8208 19372
rect 7975 19332 8208 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 7248 19320 7254 19323
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 3568 19264 6408 19292
rect 6656 19264 7512 19292
rect 3568 19252 3574 19264
rect 6380 19156 6408 19264
rect 7374 19184 7380 19236
rect 7432 19184 7438 19236
rect 7484 19233 7512 19264
rect 8110 19252 8116 19304
rect 8168 19252 8174 19304
rect 8312 19292 8340 19400
rect 8754 19388 8760 19440
rect 8812 19428 8818 19440
rect 10045 19431 10103 19437
rect 8812 19400 9536 19428
rect 8812 19388 8818 19400
rect 9508 19369 9536 19400
rect 10045 19397 10057 19431
rect 10091 19428 10103 19431
rect 10428 19428 10456 19468
rect 10091 19400 10456 19428
rect 10091 19397 10103 19400
rect 10045 19391 10103 19397
rect 10962 19388 10968 19440
rect 11020 19428 11026 19440
rect 11149 19431 11207 19437
rect 11149 19428 11161 19431
rect 11020 19400 11161 19428
rect 11020 19388 11026 19400
rect 11149 19397 11161 19400
rect 11195 19397 11207 19431
rect 11256 19428 11284 19468
rect 11514 19456 11520 19508
rect 11572 19456 11578 19508
rect 12250 19456 12256 19508
rect 12308 19456 12314 19508
rect 13538 19456 13544 19508
rect 13596 19496 13602 19508
rect 14185 19499 14243 19505
rect 14185 19496 14197 19499
rect 13596 19468 14197 19496
rect 13596 19456 13602 19468
rect 14185 19465 14197 19468
rect 14231 19465 14243 19499
rect 14185 19459 14243 19465
rect 14274 19456 14280 19508
rect 14332 19496 14338 19508
rect 14553 19499 14611 19505
rect 14553 19496 14565 19499
rect 14332 19468 14565 19496
rect 14332 19456 14338 19468
rect 14553 19465 14565 19468
rect 14599 19465 14611 19499
rect 14553 19459 14611 19465
rect 14642 19456 14648 19508
rect 14700 19456 14706 19508
rect 18046 19456 18052 19508
rect 18104 19496 18110 19508
rect 18601 19499 18659 19505
rect 18601 19496 18613 19499
rect 18104 19468 18613 19496
rect 18104 19456 18110 19468
rect 18601 19465 18613 19468
rect 18647 19465 18659 19499
rect 18601 19459 18659 19465
rect 20162 19456 20168 19508
rect 20220 19496 20226 19508
rect 20457 19499 20515 19505
rect 20457 19496 20469 19499
rect 20220 19468 20469 19496
rect 20220 19456 20226 19468
rect 20457 19465 20469 19468
rect 20503 19465 20515 19499
rect 20457 19459 20515 19465
rect 20625 19499 20683 19505
rect 20625 19465 20637 19499
rect 20671 19496 20683 19499
rect 21174 19496 21180 19508
rect 20671 19468 21180 19496
rect 20671 19465 20683 19468
rect 20625 19459 20683 19465
rect 21174 19456 21180 19468
rect 21232 19456 21238 19508
rect 21821 19499 21879 19505
rect 21821 19465 21833 19499
rect 21867 19496 21879 19499
rect 22462 19496 22468 19508
rect 21867 19468 22468 19496
rect 21867 19465 21879 19468
rect 21821 19459 21879 19465
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 12268 19428 12296 19456
rect 11256 19400 12296 19428
rect 12980 19431 13038 19437
rect 11149 19391 11207 19397
rect 12980 19397 12992 19431
rect 13026 19428 13038 19431
rect 13078 19428 13084 19440
rect 13026 19400 13084 19428
rect 13026 19397 13038 19400
rect 12980 19391 13038 19397
rect 13078 19388 13084 19400
rect 13136 19388 13142 19440
rect 14090 19388 14096 19440
rect 14148 19428 14154 19440
rect 14148 19400 15976 19428
rect 14148 19388 14154 19400
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 9950 19320 9956 19372
rect 10008 19320 10014 19372
rect 10410 19320 10416 19372
rect 10468 19320 10474 19372
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 11747 19332 11836 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8312 19264 9045 19292
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 9140 19264 10180 19292
rect 7469 19227 7527 19233
rect 7469 19193 7481 19227
rect 7515 19193 7527 19227
rect 7469 19187 7527 19193
rect 7558 19184 7564 19236
rect 7616 19224 7622 19236
rect 8128 19224 8156 19252
rect 9140 19224 9168 19264
rect 7616 19196 8156 19224
rect 8220 19196 9168 19224
rect 9217 19227 9275 19233
rect 7616 19184 7622 19196
rect 8220 19156 8248 19196
rect 9217 19193 9229 19227
rect 9263 19224 9275 19227
rect 9674 19224 9680 19236
rect 9263 19196 9680 19224
rect 9263 19193 9275 19196
rect 9217 19187 9275 19193
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 10152 19224 10180 19264
rect 10226 19252 10232 19304
rect 10284 19292 10290 19304
rect 10686 19292 10692 19304
rect 10284 19264 10692 19292
rect 10284 19252 10290 19264
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 11422 19224 11428 19236
rect 10152 19196 11428 19224
rect 11422 19184 11428 19196
rect 11480 19184 11486 19236
rect 11808 19233 11836 19332
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12158 19360 12164 19372
rect 11940 19332 12164 19360
rect 11940 19320 11946 19332
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12713 19363 12771 19369
rect 12713 19360 12725 19363
rect 12584 19332 12725 19360
rect 12584 19320 12590 19332
rect 12713 19329 12725 19332
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 15948 19369 15976 19400
rect 16758 19388 16764 19440
rect 16816 19388 16822 19440
rect 18414 19428 18420 19440
rect 17236 19400 18420 19428
rect 15933 19363 15991 19369
rect 14056 19332 14136 19360
rect 14056 19320 14062 19332
rect 12345 19295 12403 19301
rect 12345 19261 12357 19295
rect 12391 19261 12403 19295
rect 12345 19255 12403 19261
rect 11793 19227 11851 19233
rect 11793 19193 11805 19227
rect 11839 19193 11851 19227
rect 11793 19187 11851 19193
rect 6380 19128 8248 19156
rect 8754 19116 8760 19168
rect 8812 19116 8818 19168
rect 9122 19116 9128 19168
rect 9180 19116 9186 19168
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9585 19159 9643 19165
rect 9585 19156 9597 19159
rect 9364 19128 9597 19156
rect 9364 19116 9370 19128
rect 9585 19125 9597 19128
rect 9631 19125 9643 19159
rect 12360 19156 12388 19255
rect 14108 19233 14136 19332
rect 15933 19329 15945 19363
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 16942 19360 16948 19372
rect 16899 19332 16948 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 17236 19369 17264 19400
rect 18414 19388 18420 19400
rect 18472 19388 18478 19440
rect 20257 19431 20315 19437
rect 20257 19397 20269 19431
rect 20303 19397 20315 19431
rect 20257 19391 20315 19397
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17359 19332 17724 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 14737 19295 14795 19301
rect 14737 19261 14749 19295
rect 14783 19261 14795 19295
rect 17696 19292 17724 19332
rect 17770 19320 17776 19372
rect 17828 19320 17834 19372
rect 18325 19363 18383 19369
rect 18325 19360 18337 19363
rect 17926 19332 18337 19360
rect 17926 19292 17954 19332
rect 18325 19329 18337 19332
rect 18371 19360 18383 19363
rect 18598 19360 18604 19372
rect 18371 19332 18604 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 18966 19320 18972 19372
rect 19024 19320 19030 19372
rect 19518 19320 19524 19372
rect 19576 19320 19582 19372
rect 19702 19320 19708 19372
rect 19760 19360 19766 19372
rect 20070 19360 20076 19372
rect 19760 19332 20076 19360
rect 19760 19320 19766 19332
rect 20070 19320 20076 19332
rect 20128 19360 20134 19372
rect 20272 19360 20300 19391
rect 20128 19332 20300 19360
rect 20128 19320 20134 19332
rect 20346 19320 20352 19372
rect 20404 19320 20410 19372
rect 22186 19320 22192 19372
rect 22244 19320 22250 19372
rect 17696 19264 17954 19292
rect 14737 19255 14795 19261
rect 14093 19227 14151 19233
rect 14093 19193 14105 19227
rect 14139 19193 14151 19227
rect 14093 19187 14151 19193
rect 14274 19156 14280 19168
rect 12360 19128 14280 19156
rect 9585 19119 9643 19125
rect 14274 19116 14280 19128
rect 14332 19156 14338 19168
rect 14752 19156 14780 19255
rect 20162 19252 20168 19304
rect 20220 19292 20226 19304
rect 20364 19292 20392 19320
rect 20220 19264 20392 19292
rect 20220 19252 20226 19264
rect 22646 19252 22652 19304
rect 22704 19292 22710 19304
rect 23293 19295 23351 19301
rect 23293 19292 23305 19295
rect 22704 19264 23305 19292
rect 22704 19252 22710 19264
rect 23293 19261 23305 19264
rect 23339 19261 23351 19295
rect 23293 19255 23351 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19261 23627 19295
rect 23569 19255 23627 19261
rect 14332 19128 14780 19156
rect 14332 19116 14338 19128
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 20441 19159 20499 19165
rect 20441 19156 20453 19159
rect 19576 19128 20453 19156
rect 19576 19116 19582 19128
rect 20441 19125 20453 19128
rect 20487 19125 20499 19159
rect 20441 19119 20499 19125
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 23584 19156 23612 19255
rect 22152 19128 23612 19156
rect 22152 19116 22158 19128
rect 1104 19066 26864 19088
rect 1104 19014 2918 19066
rect 2970 19014 2982 19066
rect 3034 19014 3046 19066
rect 3098 19014 3110 19066
rect 3162 19014 3174 19066
rect 3226 19014 3238 19066
rect 3290 19014 6918 19066
rect 6970 19014 6982 19066
rect 7034 19014 7046 19066
rect 7098 19014 7110 19066
rect 7162 19014 7174 19066
rect 7226 19014 7238 19066
rect 7290 19014 10918 19066
rect 10970 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 11238 19066
rect 11290 19014 14918 19066
rect 14970 19014 14982 19066
rect 15034 19014 15046 19066
rect 15098 19014 15110 19066
rect 15162 19014 15174 19066
rect 15226 19014 15238 19066
rect 15290 19014 18918 19066
rect 18970 19014 18982 19066
rect 19034 19014 19046 19066
rect 19098 19014 19110 19066
rect 19162 19014 19174 19066
rect 19226 19014 19238 19066
rect 19290 19014 22918 19066
rect 22970 19014 22982 19066
rect 23034 19014 23046 19066
rect 23098 19014 23110 19066
rect 23162 19014 23174 19066
rect 23226 19014 23238 19066
rect 23290 19014 26864 19066
rect 1104 18992 26864 19014
rect 4982 18912 4988 18964
rect 5040 18952 5046 18964
rect 8481 18955 8539 18961
rect 5040 18924 8064 18952
rect 5040 18912 5046 18924
rect 8036 18884 8064 18924
rect 8481 18921 8493 18955
rect 8527 18952 8539 18955
rect 9122 18952 9128 18964
rect 8527 18924 9128 18952
rect 8527 18921 8539 18924
rect 8481 18915 8539 18921
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 9858 18952 9864 18964
rect 9692 18924 9864 18952
rect 9692 18884 9720 18924
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 9950 18912 9956 18964
rect 10008 18952 10014 18964
rect 10778 18952 10784 18964
rect 10008 18924 10784 18952
rect 10008 18912 10014 18924
rect 10778 18912 10784 18924
rect 10836 18952 10842 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10836 18924 11069 18952
rect 10836 18912 10842 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 12066 18912 12072 18964
rect 12124 18952 12130 18964
rect 12161 18955 12219 18961
rect 12161 18952 12173 18955
rect 12124 18924 12173 18952
rect 12124 18912 12130 18924
rect 12161 18921 12173 18924
rect 12207 18921 12219 18955
rect 17034 18952 17040 18964
rect 12161 18915 12219 18921
rect 12406 18924 17040 18952
rect 8036 18856 9720 18884
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 5074 18816 5080 18828
rect 4663 18788 5080 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 6546 18776 6552 18828
rect 6604 18816 6610 18828
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 6604 18788 7573 18816
rect 6604 18776 6610 18788
rect 7561 18785 7573 18788
rect 7607 18785 7619 18819
rect 7561 18779 7619 18785
rect 7760 18788 7972 18816
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18748 2375 18751
rect 3510 18748 3516 18760
rect 2363 18720 3516 18748
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 3510 18708 3516 18720
rect 3568 18708 3574 18760
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18748 3663 18751
rect 3651 18720 4016 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 2130 18572 2136 18624
rect 2188 18572 2194 18624
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 3988 18621 4016 18720
rect 4798 18708 4804 18760
rect 4856 18708 4862 18760
rect 4890 18708 4896 18760
rect 4948 18708 4954 18760
rect 5258 18708 5264 18760
rect 5316 18757 5322 18760
rect 5316 18748 5324 18757
rect 6917 18751 6975 18757
rect 5316 18720 5361 18748
rect 5316 18711 5324 18720
rect 6917 18717 6929 18751
rect 6963 18748 6975 18751
rect 7190 18748 7196 18760
rect 6963 18720 7196 18748
rect 6963 18717 6975 18720
rect 6917 18711 6975 18717
rect 5316 18708 5322 18711
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18748 7435 18751
rect 7466 18748 7472 18760
rect 7423 18720 7472 18748
rect 7423 18717 7435 18720
rect 7377 18711 7435 18717
rect 7466 18708 7472 18720
rect 7524 18748 7530 18760
rect 7760 18748 7788 18788
rect 7944 18757 7972 18788
rect 7524 18720 7788 18748
rect 7837 18751 7895 18757
rect 7524 18708 7530 18720
rect 7837 18717 7849 18751
rect 7883 18717 7895 18751
rect 7837 18711 7895 18717
rect 7930 18751 7988 18757
rect 7930 18717 7942 18751
rect 7976 18717 7988 18751
rect 8036 18748 8064 18856
rect 10686 18844 10692 18896
rect 10744 18884 10750 18896
rect 12406 18884 12434 18924
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 22186 18912 22192 18964
rect 22244 18912 22250 18964
rect 26418 18912 26424 18964
rect 26476 18912 26482 18964
rect 10744 18856 12434 18884
rect 10744 18844 10750 18856
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 8812 18788 9812 18816
rect 8812 18776 8818 18788
rect 8113 18751 8171 18757
rect 8113 18748 8125 18751
rect 8036 18720 8125 18748
rect 7930 18711 7988 18717
rect 8113 18717 8125 18720
rect 8159 18717 8171 18751
rect 8113 18711 8171 18717
rect 8343 18751 8401 18757
rect 8343 18717 8355 18751
rect 8389 18748 8401 18751
rect 8478 18748 8484 18760
rect 8389 18720 8484 18748
rect 8389 18717 8401 18720
rect 8343 18711 8401 18717
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 4396 18652 4568 18680
rect 4396 18640 4402 18652
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 2832 18584 3433 18612
rect 2832 18572 2838 18584
rect 3421 18581 3433 18584
rect 3467 18581 3479 18615
rect 3421 18575 3479 18581
rect 3973 18615 4031 18621
rect 3973 18581 3985 18615
rect 4019 18581 4031 18615
rect 3973 18575 4031 18581
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 4433 18615 4491 18621
rect 4433 18612 4445 18615
rect 4304 18584 4445 18612
rect 4304 18572 4310 18584
rect 4433 18581 4445 18584
rect 4479 18581 4491 18615
rect 4540 18612 4568 18652
rect 4982 18640 4988 18692
rect 5040 18680 5046 18692
rect 5077 18683 5135 18689
rect 5077 18680 5089 18683
rect 5040 18652 5089 18680
rect 5040 18640 5046 18652
rect 5077 18649 5089 18652
rect 5123 18649 5135 18683
rect 5077 18643 5135 18649
rect 5169 18683 5227 18689
rect 5169 18649 5181 18683
rect 5215 18649 5227 18683
rect 5169 18643 5227 18649
rect 5184 18612 5212 18643
rect 7558 18640 7564 18692
rect 7616 18680 7622 18692
rect 7852 18680 7880 18711
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 9033 18751 9091 18757
rect 9033 18717 9045 18751
rect 9079 18748 9091 18751
rect 9306 18748 9312 18760
rect 9079 18720 9312 18748
rect 9079 18717 9091 18720
rect 9033 18711 9091 18717
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 9674 18708 9680 18760
rect 9732 18708 9738 18760
rect 9784 18748 9812 18788
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14737 18819 14795 18825
rect 14737 18816 14749 18819
rect 14148 18788 14749 18816
rect 14148 18776 14154 18788
rect 14737 18785 14749 18788
rect 14783 18785 14795 18819
rect 14737 18779 14795 18785
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 9784 18720 11621 18748
rect 11609 18717 11621 18720
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 11701 18751 11759 18757
rect 11701 18717 11713 18751
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 7616 18652 7880 18680
rect 7616 18640 7622 18652
rect 8202 18640 8208 18692
rect 8260 18640 8266 18692
rect 8496 18680 8524 18708
rect 9122 18680 9128 18692
rect 8496 18652 9128 18680
rect 9122 18640 9128 18652
rect 9180 18640 9186 18692
rect 9922 18683 9980 18689
rect 9922 18680 9934 18683
rect 9232 18652 9934 18680
rect 4540 18584 5212 18612
rect 5445 18615 5503 18621
rect 4433 18575 4491 18581
rect 5445 18581 5457 18615
rect 5491 18612 5503 18615
rect 5534 18612 5540 18624
rect 5491 18584 5540 18612
rect 5491 18581 5503 18584
rect 5445 18575 5503 18581
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 6733 18615 6791 18621
rect 6733 18581 6745 18615
rect 6779 18612 6791 18615
rect 6914 18612 6920 18624
rect 6779 18584 6920 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7006 18572 7012 18624
rect 7064 18572 7070 18624
rect 7469 18615 7527 18621
rect 7469 18581 7481 18615
rect 7515 18612 7527 18615
rect 8294 18612 8300 18624
rect 7515 18584 8300 18612
rect 7515 18581 7527 18584
rect 7469 18575 7527 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 9232 18621 9260 18652
rect 9922 18649 9934 18652
rect 9968 18649 9980 18683
rect 11716 18680 11744 18711
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18748 12035 18751
rect 12066 18748 12072 18760
rect 12023 18720 12072 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12066 18708 12072 18720
rect 12124 18748 12130 18760
rect 14366 18748 14372 18760
rect 12124 18720 14372 18748
rect 12124 18708 12130 18720
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14752 18748 14780 18779
rect 17586 18776 17592 18828
rect 17644 18776 17650 18828
rect 18138 18816 18144 18828
rect 18064 18788 18144 18816
rect 18064 18757 18092 18788
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19392 18788 19441 18816
rect 19392 18776 19398 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 19429 18779 19487 18785
rect 16577 18751 16635 18757
rect 16577 18748 16589 18751
rect 14752 18720 16589 18748
rect 16577 18717 16589 18720
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18598 18708 18604 18760
rect 18656 18748 18662 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18656 18720 19257 18748
rect 18656 18708 18662 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 22097 18751 22155 18757
rect 22097 18717 22109 18751
rect 22143 18748 22155 18751
rect 22554 18748 22560 18760
rect 22143 18720 22560 18748
rect 22143 18717 22155 18720
rect 22097 18711 22155 18717
rect 22554 18708 22560 18720
rect 22612 18708 22618 18760
rect 23382 18708 23388 18760
rect 23440 18748 23446 18760
rect 24673 18751 24731 18757
rect 24673 18748 24685 18751
rect 23440 18720 24685 18748
rect 23440 18708 23446 18720
rect 24673 18717 24685 18720
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 12986 18680 12992 18692
rect 11716 18652 12992 18680
rect 9922 18643 9980 18649
rect 12986 18640 12992 18652
rect 13044 18640 13050 18692
rect 15004 18683 15062 18689
rect 15004 18649 15016 18683
rect 15050 18680 15062 18683
rect 15102 18680 15108 18692
rect 15050 18652 15108 18680
rect 15050 18649 15062 18652
rect 15004 18643 15062 18649
rect 15102 18640 15108 18652
rect 15160 18640 15166 18692
rect 17405 18683 17463 18689
rect 17405 18649 17417 18683
rect 17451 18680 17463 18683
rect 17494 18680 17500 18692
rect 17451 18652 17500 18680
rect 17451 18649 17463 18652
rect 17405 18643 17463 18649
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 17678 18640 17684 18692
rect 17736 18640 17742 18692
rect 18141 18683 18199 18689
rect 18141 18649 18153 18683
rect 18187 18649 18199 18683
rect 18141 18643 18199 18649
rect 18233 18683 18291 18689
rect 18233 18649 18245 18683
rect 18279 18680 18291 18683
rect 18690 18680 18696 18692
rect 18279 18652 18696 18680
rect 18279 18649 18291 18652
rect 18233 18643 18291 18649
rect 9217 18615 9275 18621
rect 9217 18581 9229 18615
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 9306 18572 9312 18624
rect 9364 18572 9370 18624
rect 16117 18615 16175 18621
rect 16117 18581 16129 18615
rect 16163 18612 16175 18615
rect 16850 18612 16856 18624
rect 16163 18584 16856 18612
rect 16163 18581 16175 18584
rect 16117 18575 16175 18581
rect 16850 18572 16856 18584
rect 16908 18572 16914 18624
rect 18156 18612 18184 18643
rect 18690 18640 18696 18652
rect 18748 18680 18754 18692
rect 18874 18680 18880 18692
rect 18748 18652 18880 18680
rect 18748 18640 18754 18652
rect 18874 18640 18880 18652
rect 18932 18640 18938 18692
rect 24949 18683 25007 18689
rect 24949 18649 24961 18683
rect 24995 18680 25007 18683
rect 25038 18680 25044 18692
rect 24995 18652 25044 18680
rect 24995 18649 25007 18652
rect 24949 18643 25007 18649
rect 25038 18640 25044 18652
rect 25096 18640 25102 18692
rect 26234 18680 26240 18692
rect 26174 18652 26240 18680
rect 26234 18640 26240 18652
rect 26292 18640 26298 18692
rect 19702 18612 19708 18624
rect 18156 18584 19708 18612
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 1104 18522 26864 18544
rect 1104 18470 3658 18522
rect 3710 18470 3722 18522
rect 3774 18470 3786 18522
rect 3838 18470 3850 18522
rect 3902 18470 3914 18522
rect 3966 18470 3978 18522
rect 4030 18470 7658 18522
rect 7710 18470 7722 18522
rect 7774 18470 7786 18522
rect 7838 18470 7850 18522
rect 7902 18470 7914 18522
rect 7966 18470 7978 18522
rect 8030 18470 11658 18522
rect 11710 18470 11722 18522
rect 11774 18470 11786 18522
rect 11838 18470 11850 18522
rect 11902 18470 11914 18522
rect 11966 18470 11978 18522
rect 12030 18470 15658 18522
rect 15710 18470 15722 18522
rect 15774 18470 15786 18522
rect 15838 18470 15850 18522
rect 15902 18470 15914 18522
rect 15966 18470 15978 18522
rect 16030 18470 19658 18522
rect 19710 18470 19722 18522
rect 19774 18470 19786 18522
rect 19838 18470 19850 18522
rect 19902 18470 19914 18522
rect 19966 18470 19978 18522
rect 20030 18470 23658 18522
rect 23710 18470 23722 18522
rect 23774 18470 23786 18522
rect 23838 18470 23850 18522
rect 23902 18470 23914 18522
rect 23966 18470 23978 18522
rect 24030 18470 26864 18522
rect 1104 18448 26864 18470
rect 3881 18411 3939 18417
rect 3881 18377 3893 18411
rect 3927 18408 3939 18411
rect 4338 18408 4344 18420
rect 3927 18380 4344 18408
rect 3927 18377 3939 18380
rect 3881 18371 3939 18377
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 5350 18368 5356 18420
rect 5408 18368 5414 18420
rect 5445 18411 5503 18417
rect 5445 18377 5457 18411
rect 5491 18377 5503 18411
rect 7006 18408 7012 18420
rect 5445 18371 5503 18377
rect 6012 18380 7012 18408
rect 4240 18343 4298 18349
rect 2516 18312 4016 18340
rect 2516 18284 2544 18312
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18272 2099 18275
rect 2225 18275 2283 18281
rect 2225 18272 2237 18275
rect 2087 18244 2237 18272
rect 2087 18241 2099 18244
rect 2041 18235 2099 18241
rect 2225 18241 2237 18244
rect 2271 18241 2283 18275
rect 2225 18235 2283 18241
rect 2498 18232 2504 18284
rect 2556 18232 2562 18284
rect 2774 18281 2780 18284
rect 2768 18235 2780 18281
rect 2832 18272 2838 18284
rect 3988 18281 4016 18312
rect 4240 18309 4252 18343
rect 4286 18340 4298 18343
rect 5460 18340 5488 18371
rect 4286 18312 5488 18340
rect 4286 18309 4298 18312
rect 4240 18303 4298 18309
rect 3973 18275 4031 18281
rect 2832 18244 2868 18272
rect 2774 18232 2780 18235
rect 2832 18232 2838 18244
rect 3973 18241 3985 18275
rect 4019 18272 4031 18275
rect 4062 18272 4068 18284
rect 4019 18244 4068 18272
rect 4019 18241 4031 18244
rect 3973 18235 4031 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 5626 18232 5632 18284
rect 5684 18232 5690 18284
rect 6012 18281 6040 18380
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7837 18411 7895 18417
rect 7837 18408 7849 18411
rect 7524 18380 7849 18408
rect 7524 18368 7530 18380
rect 7837 18377 7849 18380
rect 7883 18377 7895 18411
rect 7837 18371 7895 18377
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 8389 18411 8447 18417
rect 8389 18408 8401 18411
rect 8352 18380 8401 18408
rect 8352 18368 8358 18380
rect 8389 18377 8401 18380
rect 8435 18377 8447 18411
rect 8389 18371 8447 18377
rect 8956 18380 9352 18408
rect 8956 18340 8984 18380
rect 6472 18312 8984 18340
rect 6472 18281 6500 18312
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 6457 18275 6515 18281
rect 6457 18241 6469 18275
rect 6503 18241 6515 18275
rect 6713 18275 6771 18281
rect 6713 18272 6725 18275
rect 6457 18235 6515 18241
rect 6564 18244 6725 18272
rect 1394 18164 1400 18216
rect 1452 18164 1458 18216
rect 6564 18204 6592 18244
rect 6713 18241 6725 18244
rect 6759 18241 6771 18275
rect 6713 18235 6771 18241
rect 7098 18232 7104 18284
rect 7156 18272 7162 18284
rect 7156 18244 7972 18272
rect 7156 18232 7162 18244
rect 6196 18176 6592 18204
rect 6196 18145 6224 18176
rect 6181 18139 6239 18145
rect 6181 18105 6193 18139
rect 6227 18105 6239 18139
rect 7944 18136 7972 18244
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8202 18272 8208 18284
rect 8076 18244 8208 18272
rect 8076 18232 8082 18244
rect 8202 18232 8208 18244
rect 8260 18272 8266 18284
rect 8956 18281 8984 18312
rect 9205 18300 9211 18352
rect 9263 18300 9269 18352
rect 9324 18340 9352 18380
rect 9766 18368 9772 18420
rect 9824 18408 9830 18420
rect 10321 18411 10379 18417
rect 10321 18408 10333 18411
rect 9824 18380 10333 18408
rect 9824 18368 9830 18380
rect 10321 18377 10333 18380
rect 10367 18377 10379 18411
rect 10321 18371 10379 18377
rect 15102 18368 15108 18420
rect 15160 18368 15166 18420
rect 15749 18411 15807 18417
rect 15749 18377 15761 18411
rect 15795 18377 15807 18411
rect 23382 18408 23388 18420
rect 15749 18371 15807 18377
rect 22204 18380 23388 18408
rect 9674 18340 9680 18352
rect 9324 18312 9680 18340
rect 9674 18300 9680 18312
rect 9732 18340 9738 18352
rect 11149 18343 11207 18349
rect 11149 18340 11161 18343
rect 9732 18312 11161 18340
rect 9732 18300 9738 18312
rect 11149 18309 11161 18312
rect 11195 18309 11207 18343
rect 11149 18303 11207 18309
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 8260 18244 8309 18272
rect 8260 18232 8266 18244
rect 8297 18241 8309 18244
rect 8343 18241 8355 18275
rect 8297 18235 8355 18241
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 9048 18244 10364 18272
rect 8570 18164 8576 18216
rect 8628 18164 8634 18216
rect 9048 18204 9076 18244
rect 8956 18176 9076 18204
rect 10336 18204 10364 18244
rect 10410 18232 10416 18284
rect 10468 18232 10474 18284
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18272 15347 18275
rect 15764 18272 15792 18371
rect 16390 18340 16396 18352
rect 15335 18244 15792 18272
rect 16040 18312 16396 18340
rect 15335 18241 15347 18244
rect 15289 18235 15347 18241
rect 12066 18204 12072 18216
rect 10336 18176 12072 18204
rect 8956 18136 8984 18176
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 14734 18164 14740 18216
rect 14792 18204 14798 18216
rect 16040 18204 16068 18312
rect 16390 18300 16396 18312
rect 16448 18300 16454 18352
rect 18138 18300 18144 18352
rect 18196 18340 18202 18352
rect 18325 18343 18383 18349
rect 18325 18340 18337 18343
rect 18196 18312 18337 18340
rect 18196 18300 18202 18312
rect 18325 18309 18337 18312
rect 18371 18309 18383 18343
rect 18325 18303 18383 18309
rect 18874 18300 18880 18352
rect 18932 18300 18938 18352
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16850 18272 16856 18284
rect 16163 18244 16856 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 17586 18232 17592 18284
rect 17644 18232 17650 18284
rect 18233 18275 18291 18281
rect 18233 18241 18245 18275
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 14792 18176 16221 18204
rect 14792 18164 14798 18176
rect 16209 18173 16221 18176
rect 16255 18173 16267 18207
rect 16209 18167 16267 18173
rect 16390 18164 16396 18216
rect 16448 18164 16454 18216
rect 16758 18164 16764 18216
rect 16816 18164 16822 18216
rect 18248 18204 18276 18235
rect 18414 18232 18420 18284
rect 18472 18232 18478 18284
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22204 18281 22232 18380
rect 23382 18368 23388 18380
rect 23440 18408 23446 18420
rect 23440 18380 24072 18408
rect 23440 18368 23446 18380
rect 23842 18340 23848 18352
rect 23690 18312 23848 18340
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 24044 18281 24072 18380
rect 25774 18368 25780 18420
rect 25832 18368 25838 18420
rect 26234 18368 26240 18420
rect 26292 18368 26298 18420
rect 24854 18300 24860 18352
rect 24912 18300 24918 18352
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 22152 18244 22201 18272
rect 22152 18232 22158 18244
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 24029 18275 24087 18281
rect 24029 18241 24041 18275
rect 24075 18241 24087 18275
rect 24029 18235 24087 18241
rect 26050 18232 26056 18284
rect 26108 18272 26114 18284
rect 26145 18275 26203 18281
rect 26145 18272 26157 18275
rect 26108 18244 26157 18272
rect 26108 18232 26114 18244
rect 26145 18241 26157 18244
rect 26191 18241 26203 18275
rect 26145 18235 26203 18241
rect 18598 18204 18604 18216
rect 18248 18176 18604 18204
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 18785 18207 18843 18213
rect 18785 18173 18797 18207
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 14826 18136 14832 18148
rect 7944 18108 8984 18136
rect 9876 18108 14832 18136
rect 6181 18099 6239 18105
rect 2317 18071 2375 18077
rect 2317 18037 2329 18071
rect 2363 18068 2375 18071
rect 4154 18068 4160 18080
rect 2363 18040 4160 18068
rect 2363 18037 2375 18040
rect 2317 18031 2375 18037
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 5166 18028 5172 18080
rect 5224 18068 5230 18080
rect 7098 18068 7104 18080
rect 5224 18040 7104 18068
rect 5224 18028 5230 18040
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7190 18028 7196 18080
rect 7248 18068 7254 18080
rect 7929 18071 7987 18077
rect 7929 18068 7941 18071
rect 7248 18040 7941 18068
rect 7248 18028 7254 18040
rect 7929 18037 7941 18040
rect 7975 18037 7987 18071
rect 7929 18031 7987 18037
rect 8110 18028 8116 18080
rect 8168 18068 8174 18080
rect 9876 18068 9904 18108
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 16114 18096 16120 18148
rect 16172 18136 16178 18148
rect 16408 18136 16436 18164
rect 16172 18108 16436 18136
rect 16172 18096 16178 18108
rect 17034 18096 17040 18148
rect 17092 18136 17098 18148
rect 17770 18136 17776 18148
rect 17092 18108 17776 18136
rect 17092 18096 17098 18108
rect 17770 18096 17776 18108
rect 17828 18096 17834 18148
rect 18138 18096 18144 18148
rect 18196 18136 18202 18148
rect 18800 18136 18828 18167
rect 22462 18164 22468 18216
rect 22520 18164 22526 18216
rect 23474 18164 23480 18216
rect 23532 18204 23538 18216
rect 24305 18207 24363 18213
rect 24305 18204 24317 18207
rect 23532 18176 24317 18204
rect 23532 18164 23538 18176
rect 24305 18173 24317 18176
rect 24351 18173 24363 18207
rect 24305 18167 24363 18173
rect 18196 18108 18828 18136
rect 18196 18096 18202 18108
rect 8168 18040 9904 18068
rect 8168 18028 8174 18040
rect 9950 18028 9956 18080
rect 10008 18068 10014 18080
rect 15378 18068 15384 18080
rect 10008 18040 15384 18068
rect 10008 18028 10014 18040
rect 15378 18028 15384 18040
rect 15436 18068 15442 18080
rect 17862 18068 17868 18080
rect 15436 18040 17868 18068
rect 15436 18028 15442 18040
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 23937 18071 23995 18077
rect 23937 18037 23949 18071
rect 23983 18068 23995 18071
rect 24118 18068 24124 18080
rect 23983 18040 24124 18068
rect 23983 18037 23995 18040
rect 23937 18031 23995 18037
rect 24118 18028 24124 18040
rect 24176 18028 24182 18080
rect 25958 18028 25964 18080
rect 26016 18028 26022 18080
rect 1104 17978 26864 18000
rect 1104 17926 2918 17978
rect 2970 17926 2982 17978
rect 3034 17926 3046 17978
rect 3098 17926 3110 17978
rect 3162 17926 3174 17978
rect 3226 17926 3238 17978
rect 3290 17926 6918 17978
rect 6970 17926 6982 17978
rect 7034 17926 7046 17978
rect 7098 17926 7110 17978
rect 7162 17926 7174 17978
rect 7226 17926 7238 17978
rect 7290 17926 10918 17978
rect 10970 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 11238 17978
rect 11290 17926 14918 17978
rect 14970 17926 14982 17978
rect 15034 17926 15046 17978
rect 15098 17926 15110 17978
rect 15162 17926 15174 17978
rect 15226 17926 15238 17978
rect 15290 17926 18918 17978
rect 18970 17926 18982 17978
rect 19034 17926 19046 17978
rect 19098 17926 19110 17978
rect 19162 17926 19174 17978
rect 19226 17926 19238 17978
rect 19290 17926 22918 17978
rect 22970 17926 22982 17978
rect 23034 17926 23046 17978
rect 23098 17926 23110 17978
rect 23162 17926 23174 17978
rect 23226 17926 23238 17978
rect 23290 17926 26864 17978
rect 1104 17904 26864 17926
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3568 17836 3801 17864
rect 3568 17824 3574 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 3789 17827 3847 17833
rect 5353 17867 5411 17873
rect 5353 17833 5365 17867
rect 5399 17864 5411 17867
rect 5626 17864 5632 17876
rect 5399 17836 5632 17864
rect 5399 17833 5411 17836
rect 5353 17827 5411 17833
rect 5626 17824 5632 17836
rect 5684 17824 5690 17876
rect 8018 17824 8024 17876
rect 8076 17824 8082 17876
rect 8570 17824 8576 17876
rect 8628 17864 8634 17876
rect 9214 17864 9220 17876
rect 8628 17836 9220 17864
rect 8628 17824 8634 17836
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 9401 17867 9459 17873
rect 9401 17833 9413 17867
rect 9447 17864 9459 17867
rect 9490 17864 9496 17876
rect 9447 17836 9496 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 10413 17867 10471 17873
rect 10413 17864 10425 17867
rect 10376 17836 10425 17864
rect 10376 17824 10382 17836
rect 10413 17833 10425 17836
rect 10459 17833 10471 17867
rect 10413 17827 10471 17833
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 17218 17864 17224 17876
rect 10652 17836 17224 17864
rect 10652 17824 10658 17836
rect 17218 17824 17224 17836
rect 17276 17864 17282 17876
rect 17678 17864 17684 17876
rect 17276 17836 17684 17864
rect 17276 17824 17282 17836
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 22094 17864 22100 17876
rect 21652 17836 22100 17864
rect 2869 17799 2927 17805
rect 2869 17765 2881 17799
rect 2915 17796 2927 17799
rect 6546 17796 6552 17808
rect 2915 17768 4200 17796
rect 2915 17765 2927 17768
rect 2869 17759 2927 17765
rect 1486 17620 1492 17672
rect 1544 17620 1550 17672
rect 1756 17663 1814 17669
rect 1756 17629 1768 17663
rect 1802 17660 1814 17663
rect 2130 17660 2136 17672
rect 1802 17632 2136 17660
rect 1802 17629 1814 17632
rect 1756 17623 1814 17629
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 4172 17669 4200 17768
rect 4356 17768 6552 17796
rect 4356 17740 4384 17768
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 11422 17756 11428 17808
rect 11480 17796 11486 17808
rect 11480 17768 12664 17796
rect 11480 17756 11486 17768
rect 4338 17688 4344 17740
rect 4396 17688 4402 17740
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17728 4859 17731
rect 4847 17700 6592 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 4890 17660 4896 17672
rect 4203 17632 4896 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17660 5043 17663
rect 5350 17660 5356 17672
rect 5031 17632 5356 17660
rect 5031 17629 5043 17632
rect 4985 17623 5043 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 4246 17552 4252 17604
rect 4304 17592 4310 17604
rect 5442 17592 5448 17604
rect 4304 17564 5448 17592
rect 4304 17552 4310 17564
rect 5442 17552 5448 17564
rect 5500 17552 5506 17604
rect 6564 17592 6592 17700
rect 6638 17688 6644 17740
rect 6696 17688 6702 17740
rect 10042 17688 10048 17740
rect 10100 17688 10106 17740
rect 10778 17688 10784 17740
rect 10836 17688 10842 17740
rect 12250 17688 12256 17740
rect 12308 17728 12314 17740
rect 12636 17737 12664 17768
rect 12437 17731 12495 17737
rect 12437 17728 12449 17731
rect 12308 17700 12449 17728
rect 12308 17688 12314 17700
rect 12437 17697 12449 17700
rect 12483 17697 12495 17731
rect 12437 17691 12495 17697
rect 12621 17731 12679 17737
rect 12621 17697 12633 17731
rect 12667 17728 12679 17731
rect 13998 17728 14004 17740
rect 12667 17700 14004 17728
rect 12667 17697 12679 17700
rect 12621 17691 12679 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 18598 17688 18604 17740
rect 18656 17688 18662 17740
rect 21652 17737 21680 17836
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 23385 17867 23443 17873
rect 23385 17833 23397 17867
rect 23431 17864 23443 17867
rect 23474 17864 23480 17876
rect 23431 17836 23480 17864
rect 23431 17833 23443 17836
rect 23385 17827 23443 17833
rect 23474 17824 23480 17836
rect 23532 17824 23538 17876
rect 23842 17824 23848 17876
rect 23900 17824 23906 17876
rect 24121 17867 24179 17873
rect 24121 17833 24133 17867
rect 24167 17864 24179 17867
rect 24854 17864 24860 17876
rect 24167 17836 24860 17864
rect 24167 17833 24179 17836
rect 24121 17827 24179 17833
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 26142 17824 26148 17876
rect 26200 17824 26206 17876
rect 21637 17731 21695 17737
rect 21637 17697 21649 17731
rect 21683 17697 21695 17731
rect 21637 17691 21695 17697
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17728 21971 17731
rect 22278 17728 22284 17740
rect 21959 17700 22284 17728
rect 21959 17697 21971 17700
rect 21913 17691 21971 17697
rect 22278 17688 22284 17700
rect 22336 17688 22342 17740
rect 22554 17688 22560 17740
rect 22612 17728 22618 17740
rect 22612 17700 23152 17728
rect 22612 17688 22618 17700
rect 6914 17669 6920 17672
rect 6908 17660 6920 17669
rect 6875 17632 6920 17660
rect 6908 17623 6920 17632
rect 6914 17620 6920 17623
rect 6972 17620 6978 17672
rect 9766 17620 9772 17672
rect 9824 17620 9830 17672
rect 10594 17620 10600 17672
rect 10652 17620 10658 17672
rect 10796 17660 10824 17688
rect 10965 17663 11023 17669
rect 10965 17660 10977 17663
rect 10796 17632 10977 17660
rect 10965 17629 10977 17632
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 13170 17660 13176 17672
rect 12391 17632 13176 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 16025 17663 16083 17669
rect 16025 17660 16037 17663
rect 14424 17632 16037 17660
rect 14424 17620 14430 17632
rect 16025 17629 16037 17632
rect 16071 17660 16083 17663
rect 16758 17660 16764 17672
rect 16071 17632 16764 17660
rect 16071 17629 16083 17632
rect 16025 17623 16083 17629
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 17954 17660 17960 17672
rect 17880 17632 17960 17660
rect 8938 17592 8944 17604
rect 6564 17564 8944 17592
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 10686 17552 10692 17604
rect 10744 17552 10750 17604
rect 10781 17595 10839 17601
rect 10781 17561 10793 17595
rect 10827 17592 10839 17595
rect 17880 17592 17908 17632
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 19242 17620 19248 17672
rect 19300 17620 19306 17672
rect 23124 17660 23152 17700
rect 23382 17688 23388 17740
rect 23440 17728 23446 17740
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 23440 17700 24409 17728
rect 23440 17688 23446 17700
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 23124 17632 23673 17660
rect 23661 17629 23673 17632
rect 23707 17660 23719 17663
rect 23937 17663 23995 17669
rect 23937 17660 23949 17663
rect 23707 17632 23949 17660
rect 23707 17629 23719 17632
rect 23661 17623 23719 17629
rect 23937 17629 23949 17632
rect 23983 17660 23995 17663
rect 24029 17663 24087 17669
rect 24029 17660 24041 17663
rect 23983 17632 24041 17660
rect 23983 17629 23995 17632
rect 23937 17623 23995 17629
rect 24029 17629 24041 17632
rect 24075 17629 24087 17663
rect 24029 17623 24087 17629
rect 10827 17564 17908 17592
rect 18325 17595 18383 17601
rect 10827 17561 10839 17564
rect 10781 17555 10839 17561
rect 18325 17561 18337 17595
rect 18371 17592 18383 17595
rect 19334 17592 19340 17604
rect 18371 17564 19340 17592
rect 18371 17561 18383 17564
rect 18325 17555 18383 17561
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 23569 17595 23627 17601
rect 23569 17592 23581 17595
rect 23138 17564 23581 17592
rect 23569 17561 23581 17564
rect 23615 17561 23627 17595
rect 23569 17555 23627 17561
rect 4798 17484 4804 17536
rect 4856 17524 4862 17536
rect 4893 17527 4951 17533
rect 4893 17524 4905 17527
rect 4856 17496 4905 17524
rect 4856 17484 4862 17496
rect 4893 17493 4905 17496
rect 4939 17493 4951 17527
rect 4893 17487 4951 17493
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 9824 17496 9873 17524
rect 9824 17484 9830 17496
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 9861 17487 9919 17493
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 11977 17527 12035 17533
rect 11977 17524 11989 17527
rect 11388 17496 11989 17524
rect 11388 17484 11394 17496
rect 11977 17493 11989 17496
rect 12023 17493 12035 17527
rect 11977 17487 12035 17493
rect 12802 17484 12808 17536
rect 12860 17524 12866 17536
rect 16114 17524 16120 17536
rect 12860 17496 16120 17524
rect 12860 17484 12866 17496
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 17957 17527 18015 17533
rect 17957 17524 17969 17527
rect 17552 17496 17969 17524
rect 17552 17484 17558 17496
rect 17957 17493 17969 17496
rect 18003 17493 18015 17527
rect 17957 17487 18015 17493
rect 18414 17484 18420 17536
rect 18472 17484 18478 17536
rect 19426 17484 19432 17536
rect 19484 17484 19490 17536
rect 24044 17524 24072 17623
rect 26050 17620 26056 17672
rect 26108 17660 26114 17672
rect 26237 17663 26295 17669
rect 26237 17660 26249 17663
rect 26108 17632 26249 17660
rect 26108 17620 26114 17632
rect 26237 17629 26249 17632
rect 26283 17629 26295 17663
rect 26237 17623 26295 17629
rect 24673 17595 24731 17601
rect 24673 17561 24685 17595
rect 24719 17592 24731 17595
rect 24762 17592 24768 17604
rect 24719 17564 24768 17592
rect 24719 17561 24731 17564
rect 24673 17555 24731 17561
rect 24762 17552 24768 17564
rect 24820 17552 24826 17604
rect 26329 17595 26387 17601
rect 26329 17592 26341 17595
rect 25898 17564 26341 17592
rect 26329 17561 26341 17564
rect 26375 17561 26387 17595
rect 26329 17555 26387 17561
rect 26050 17524 26056 17536
rect 24044 17496 26056 17524
rect 26050 17484 26056 17496
rect 26108 17484 26114 17536
rect 1104 17434 26864 17456
rect 1104 17382 3658 17434
rect 3710 17382 3722 17434
rect 3774 17382 3786 17434
rect 3838 17382 3850 17434
rect 3902 17382 3914 17434
rect 3966 17382 3978 17434
rect 4030 17382 7658 17434
rect 7710 17382 7722 17434
rect 7774 17382 7786 17434
rect 7838 17382 7850 17434
rect 7902 17382 7914 17434
rect 7966 17382 7978 17434
rect 8030 17382 11658 17434
rect 11710 17382 11722 17434
rect 11774 17382 11786 17434
rect 11838 17382 11850 17434
rect 11902 17382 11914 17434
rect 11966 17382 11978 17434
rect 12030 17382 15658 17434
rect 15710 17382 15722 17434
rect 15774 17382 15786 17434
rect 15838 17382 15850 17434
rect 15902 17382 15914 17434
rect 15966 17382 15978 17434
rect 16030 17382 19658 17434
rect 19710 17382 19722 17434
rect 19774 17382 19786 17434
rect 19838 17382 19850 17434
rect 19902 17382 19914 17434
rect 19966 17382 19978 17434
rect 20030 17382 23658 17434
rect 23710 17382 23722 17434
rect 23774 17382 23786 17434
rect 23838 17382 23850 17434
rect 23902 17382 23914 17434
rect 23966 17382 23978 17434
rect 24030 17382 26864 17434
rect 1104 17360 26864 17382
rect 3053 17323 3111 17329
rect 3053 17289 3065 17323
rect 3099 17289 3111 17323
rect 3053 17283 3111 17289
rect 1486 17212 1492 17264
rect 1544 17252 1550 17264
rect 2498 17252 2504 17264
rect 1544 17224 2504 17252
rect 1544 17212 1550 17224
rect 1688 17193 1716 17224
rect 2498 17212 2504 17224
rect 2556 17212 2562 17264
rect 3068 17252 3096 17283
rect 12986 17280 12992 17332
rect 13044 17280 13050 17332
rect 17681 17323 17739 17329
rect 17681 17289 17693 17323
rect 17727 17289 17739 17323
rect 17681 17283 17739 17289
rect 19153 17323 19211 17329
rect 19153 17289 19165 17323
rect 19199 17320 19211 17323
rect 19334 17320 19340 17332
rect 19199 17292 19340 17320
rect 19199 17289 19211 17292
rect 19153 17283 19211 17289
rect 3513 17255 3571 17261
rect 3513 17252 3525 17255
rect 3068 17224 3525 17252
rect 3513 17221 3525 17224
rect 3559 17252 3571 17255
rect 4614 17252 4620 17264
rect 3559 17224 4620 17252
rect 3559 17221 3571 17224
rect 3513 17215 3571 17221
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 6730 17212 6736 17264
rect 6788 17252 6794 17264
rect 10226 17252 10232 17264
rect 6788 17224 10232 17252
rect 6788 17212 6794 17224
rect 10226 17212 10232 17224
rect 10284 17252 10290 17264
rect 12529 17255 12587 17261
rect 10284 17224 12434 17252
rect 10284 17212 10290 17224
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 1940 17187 1998 17193
rect 1940 17153 1952 17187
rect 1986 17184 1998 17187
rect 2222 17184 2228 17196
rect 1986 17156 2228 17184
rect 1986 17153 1998 17156
rect 1940 17147 1998 17153
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4798 17184 4804 17196
rect 4212 17156 4804 17184
rect 4212 17144 4218 17156
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9732 17156 9781 17184
rect 9732 17144 9738 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 10502 17144 10508 17196
rect 10560 17144 10566 17196
rect 12406 17184 12434 17224
rect 12529 17221 12541 17255
rect 12575 17252 12587 17255
rect 17126 17252 17132 17264
rect 12575 17224 13308 17252
rect 12575 17221 12587 17224
rect 12529 17215 12587 17221
rect 13280 17196 13308 17224
rect 13372 17224 17132 17252
rect 13173 17187 13231 17193
rect 13173 17184 13185 17187
rect 12406 17156 13185 17184
rect 13173 17153 13185 17156
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 3605 17119 3663 17125
rect 3605 17116 3617 17119
rect 3436 17088 3617 17116
rect 2774 17008 2780 17060
rect 2832 17048 2838 17060
rect 3145 17051 3203 17057
rect 3145 17048 3157 17051
rect 2832 17020 3157 17048
rect 2832 17008 2838 17020
rect 3145 17017 3157 17020
rect 3191 17017 3203 17051
rect 3145 17011 3203 17017
rect 3436 16980 3464 17088
rect 3605 17085 3617 17088
rect 3651 17085 3663 17119
rect 3605 17079 3663 17085
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 4338 17116 4344 17128
rect 3743 17088 4344 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 3510 17008 3516 17060
rect 3568 17048 3574 17060
rect 3712 17048 3740 17079
rect 4338 17076 4344 17088
rect 4396 17076 4402 17128
rect 12618 17076 12624 17128
rect 12676 17076 12682 17128
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17116 12863 17119
rect 12894 17116 12900 17128
rect 12851 17088 12900 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 3568 17020 3740 17048
rect 3568 17008 3574 17020
rect 8938 17008 8944 17060
rect 8996 17048 9002 17060
rect 9490 17048 9496 17060
rect 8996 17020 9496 17048
rect 8996 17008 9002 17020
rect 9490 17008 9496 17020
rect 9548 17048 9554 17060
rect 12820 17048 12848 17079
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13188 17116 13216 17147
rect 13262 17144 13268 17196
rect 13320 17144 13326 17196
rect 13372 17116 13400 17224
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 17696 17252 17724 17283
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 21821 17323 21879 17329
rect 21821 17289 21833 17323
rect 21867 17320 21879 17323
rect 22462 17320 22468 17332
rect 21867 17292 22468 17320
rect 21867 17289 21879 17292
rect 21821 17283 21879 17289
rect 22462 17280 22468 17292
rect 22520 17280 22526 17332
rect 24581 17323 24639 17329
rect 24581 17289 24593 17323
rect 24627 17320 24639 17323
rect 25038 17320 25044 17332
rect 24627 17292 25044 17320
rect 24627 17289 24639 17292
rect 24581 17283 24639 17289
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 18018 17255 18076 17261
rect 18018 17252 18030 17255
rect 17696 17224 18030 17252
rect 18018 17221 18030 17224
rect 18064 17221 18076 17255
rect 18018 17215 18076 17221
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 20358 17255 20416 17261
rect 20358 17252 20370 17255
rect 19484 17224 20370 17252
rect 19484 17212 19490 17224
rect 20358 17221 20370 17224
rect 20404 17221 20416 17255
rect 20358 17215 20416 17221
rect 22830 17212 22836 17264
rect 22888 17212 22894 17264
rect 23293 17255 23351 17261
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 23382 17252 23388 17264
rect 23339 17224 23388 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 25958 17252 25964 17264
rect 25622 17224 25964 17252
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 13722 17184 13728 17196
rect 13587 17156 13728 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 13188 17088 13400 17116
rect 13464 17116 13492 17147
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17184 14335 17187
rect 14366 17184 14372 17196
rect 14323 17156 14372 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 14550 17193 14556 17196
rect 14544 17147 14556 17193
rect 14550 17144 14556 17147
rect 14608 17144 14614 17196
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 15672 17156 15761 17184
rect 13814 17116 13820 17128
rect 13464 17088 13820 17116
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 9548 17020 12848 17048
rect 9548 17008 9554 17020
rect 4341 16983 4399 16989
rect 4341 16980 4353 16983
rect 3436 16952 4353 16980
rect 4341 16949 4353 16952
rect 4387 16980 4399 16983
rect 4430 16980 4436 16992
rect 4387 16952 4436 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 10318 16940 10324 16992
rect 10376 16940 10382 16992
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11572 16952 12173 16980
rect 11572 16940 11578 16952
rect 12161 16949 12173 16952
rect 12207 16949 12219 16983
rect 12161 16943 12219 16949
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15672 16989 15700 17156
rect 15749 17153 15761 17156
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 15948 17116 15976 17147
rect 16022 17144 16028 17196
rect 16080 17144 16086 17196
rect 16114 17144 16120 17196
rect 16172 17144 16178 17196
rect 17494 17144 17500 17196
rect 17552 17144 17558 17196
rect 21637 17187 21695 17193
rect 21637 17153 21649 17187
rect 21683 17184 21695 17187
rect 21683 17156 22094 17184
rect 21683 17153 21695 17156
rect 21637 17147 21695 17153
rect 16482 17116 16488 17128
rect 15948 17088 16488 17116
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 17678 17116 17684 17128
rect 16816 17088 17684 17116
rect 16816 17076 16822 17088
rect 17678 17076 17684 17088
rect 17736 17116 17742 17128
rect 17773 17119 17831 17125
rect 17773 17116 17785 17119
rect 17736 17088 17785 17116
rect 17736 17076 17742 17088
rect 17773 17085 17785 17088
rect 17819 17085 17831 17119
rect 17773 17079 17831 17085
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 21542 17116 21548 17128
rect 20671 17088 21548 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 21542 17076 21548 17088
rect 21600 17076 21606 17128
rect 22066 17116 22094 17156
rect 22554 17116 22560 17128
rect 22066 17088 22560 17116
rect 22554 17076 22560 17088
rect 22612 17076 22618 17128
rect 23569 17119 23627 17125
rect 23569 17085 23581 17119
rect 23615 17085 23627 17119
rect 23569 17079 23627 17085
rect 23584 17048 23612 17079
rect 26050 17076 26056 17128
rect 26108 17076 26114 17128
rect 26329 17119 26387 17125
rect 26329 17085 26341 17119
rect 26375 17085 26387 17119
rect 26329 17079 26387 17085
rect 23584 17020 25084 17048
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15528 16952 15669 16980
rect 15528 16940 15534 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 15657 16943 15715 16949
rect 16301 16983 16359 16989
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 16666 16980 16672 16992
rect 16347 16952 16672 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 19245 16983 19303 16989
rect 19245 16949 19257 16983
rect 19291 16980 19303 16983
rect 19426 16980 19432 16992
rect 19291 16952 19432 16980
rect 19291 16949 19303 16952
rect 19245 16943 19303 16949
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 21450 16940 21456 16992
rect 21508 16980 21514 16992
rect 21545 16983 21603 16989
rect 21545 16980 21557 16983
rect 21508 16952 21557 16980
rect 21508 16940 21514 16952
rect 21545 16949 21557 16952
rect 21591 16949 21603 16983
rect 21545 16943 21603 16949
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 23584 16980 23612 17020
rect 22152 16952 23612 16980
rect 25056 16980 25084 17020
rect 26344 16980 26372 17079
rect 25056 16952 26372 16980
rect 22152 16940 22158 16952
rect 1104 16890 26864 16912
rect 1104 16838 2918 16890
rect 2970 16838 2982 16890
rect 3034 16838 3046 16890
rect 3098 16838 3110 16890
rect 3162 16838 3174 16890
rect 3226 16838 3238 16890
rect 3290 16838 6918 16890
rect 6970 16838 6982 16890
rect 7034 16838 7046 16890
rect 7098 16838 7110 16890
rect 7162 16838 7174 16890
rect 7226 16838 7238 16890
rect 7290 16838 10918 16890
rect 10970 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 11238 16890
rect 11290 16838 14918 16890
rect 14970 16838 14982 16890
rect 15034 16838 15046 16890
rect 15098 16838 15110 16890
rect 15162 16838 15174 16890
rect 15226 16838 15238 16890
rect 15290 16838 18918 16890
rect 18970 16838 18982 16890
rect 19034 16838 19046 16890
rect 19098 16838 19110 16890
rect 19162 16838 19174 16890
rect 19226 16838 19238 16890
rect 19290 16838 22918 16890
rect 22970 16838 22982 16890
rect 23034 16838 23046 16890
rect 23098 16838 23110 16890
rect 23162 16838 23174 16890
rect 23226 16838 23238 16890
rect 23290 16838 26864 16890
rect 1104 16816 26864 16838
rect 2222 16736 2228 16788
rect 2280 16736 2286 16788
rect 4893 16779 4951 16785
rect 4893 16745 4905 16779
rect 4939 16776 4951 16779
rect 5994 16776 6000 16788
rect 4939 16748 6000 16776
rect 4939 16745 4951 16748
rect 4893 16739 4951 16745
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 9732 16748 10640 16776
rect 9732 16736 9738 16748
rect 8202 16708 8208 16720
rect 6748 16680 8208 16708
rect 4982 16600 4988 16652
rect 5040 16600 5046 16652
rect 6748 16649 6776 16680
rect 8202 16668 8208 16680
rect 8260 16668 8266 16720
rect 10612 16708 10640 16748
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 10744 16748 11069 16776
rect 10744 16736 10750 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11057 16739 11115 16745
rect 13173 16779 13231 16785
rect 13173 16745 13185 16779
rect 13219 16776 13231 16779
rect 13262 16776 13268 16788
rect 13219 16748 13268 16776
rect 13219 16745 13231 16748
rect 13173 16739 13231 16745
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 13814 16736 13820 16788
rect 13872 16736 13878 16788
rect 16482 16776 16488 16788
rect 15212 16748 16488 16776
rect 10962 16708 10968 16720
rect 10612 16680 10968 16708
rect 10962 16668 10968 16680
rect 11020 16708 11026 16720
rect 15212 16708 15240 16748
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 18414 16776 18420 16788
rect 17604 16748 18420 16776
rect 11020 16680 11836 16708
rect 11020 16668 11026 16680
rect 6733 16643 6791 16649
rect 6733 16609 6745 16643
rect 6779 16609 6791 16643
rect 6733 16603 6791 16609
rect 6822 16600 6828 16652
rect 6880 16600 6886 16652
rect 9674 16600 9680 16652
rect 9732 16600 9738 16652
rect 11808 16649 11836 16680
rect 13648 16680 15240 16708
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 13648 16640 13676 16680
rect 11793 16603 11851 16609
rect 13556 16612 13676 16640
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 2774 16572 2780 16584
rect 2455 16544 2780 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 4246 16532 4252 16584
rect 4304 16532 4310 16584
rect 4338 16532 4344 16584
rect 4396 16532 4402 16584
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 4755 16575 4813 16581
rect 4755 16541 4767 16575
rect 4801 16572 4813 16575
rect 5000 16572 5028 16600
rect 5350 16572 5356 16584
rect 4801 16544 5356 16572
rect 4801 16541 4813 16544
rect 4755 16535 4813 16541
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 6641 16575 6699 16581
rect 6641 16541 6653 16575
rect 6687 16572 6699 16575
rect 7098 16572 7104 16584
rect 6687 16544 7104 16572
rect 6687 16541 6699 16544
rect 6641 16535 6699 16541
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 7469 16575 7527 16581
rect 7469 16572 7481 16575
rect 7208 16544 7481 16572
rect 4525 16507 4583 16513
rect 4525 16473 4537 16507
rect 4571 16473 4583 16507
rect 4525 16467 4583 16473
rect 4540 16436 4568 16467
rect 4982 16464 4988 16516
rect 5040 16504 5046 16516
rect 7208 16504 7236 16544
rect 7469 16541 7481 16544
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 9944 16575 10002 16581
rect 9944 16541 9956 16575
rect 9990 16572 10002 16575
rect 10318 16572 10324 16584
rect 9990 16544 10324 16572
rect 9990 16541 10002 16544
rect 9944 16535 10002 16541
rect 5040 16476 7236 16504
rect 5040 16464 5046 16476
rect 7282 16464 7288 16516
rect 7340 16464 7346 16516
rect 7374 16464 7380 16516
rect 7432 16464 7438 16516
rect 7484 16504 7512 16535
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 11241 16575 11299 16581
rect 11241 16541 11253 16575
rect 11287 16572 11299 16575
rect 11330 16572 11336 16584
rect 11287 16544 11336 16572
rect 11287 16541 11299 16544
rect 11241 16535 11299 16541
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 11514 16532 11520 16584
rect 11572 16532 11578 16584
rect 11624 16544 12296 16572
rect 11624 16504 11652 16544
rect 12268 16516 12296 16544
rect 13170 16532 13176 16584
rect 13228 16572 13234 16584
rect 13265 16575 13323 16581
rect 13265 16572 13277 16575
rect 13228 16544 13277 16572
rect 13228 16532 13234 16544
rect 13265 16541 13277 16544
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13556 16572 13584 16612
rect 14826 16600 14832 16652
rect 14884 16640 14890 16652
rect 15013 16643 15071 16649
rect 15013 16640 15025 16643
rect 14884 16612 15025 16640
rect 14884 16600 14890 16612
rect 15013 16609 15025 16612
rect 15059 16609 15071 16643
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15013 16603 15071 16609
rect 15120 16612 15301 16640
rect 13495 16544 13584 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 13630 16532 13636 16584
rect 13688 16532 13694 16584
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16541 14243 16575
rect 14185 16535 14243 16541
rect 12038 16507 12096 16513
rect 12038 16504 12050 16507
rect 7484 16476 11652 16504
rect 11716 16476 12050 16504
rect 5258 16436 5264 16448
rect 4540 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5902 16396 5908 16448
rect 5960 16436 5966 16448
rect 6273 16439 6331 16445
rect 6273 16436 6285 16439
rect 5960 16408 6285 16436
rect 5960 16396 5966 16408
rect 6273 16405 6285 16408
rect 6319 16405 6331 16439
rect 6273 16399 6331 16405
rect 7558 16396 7564 16448
rect 7616 16436 7622 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7616 16408 7665 16436
rect 7616 16396 7622 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 7653 16399 7711 16405
rect 11422 16396 11428 16448
rect 11480 16396 11486 16448
rect 11716 16445 11744 16476
rect 12038 16473 12050 16476
rect 12084 16473 12096 16507
rect 12038 16467 12096 16473
rect 12250 16464 12256 16516
rect 12308 16464 12314 16516
rect 13538 16464 13544 16516
rect 13596 16464 13602 16516
rect 14200 16504 14228 16535
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 15120 16572 15148 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 16632 16612 17325 16640
rect 16632 16600 16638 16612
rect 17313 16609 17325 16612
rect 17359 16609 17371 16643
rect 17604 16640 17632 16748
rect 18414 16736 18420 16748
rect 18472 16776 18478 16788
rect 18472 16748 18644 16776
rect 18472 16736 18478 16748
rect 18616 16708 18644 16748
rect 19242 16736 19248 16788
rect 19300 16736 19306 16788
rect 20070 16736 20076 16788
rect 20128 16736 20134 16788
rect 22094 16776 22100 16788
rect 20732 16748 22100 16776
rect 19610 16708 19616 16720
rect 18616 16680 19616 16708
rect 19610 16668 19616 16680
rect 19668 16668 19674 16720
rect 20622 16708 20628 16720
rect 19904 16680 20628 16708
rect 17313 16603 17371 16609
rect 17420 16612 17632 16640
rect 16022 16572 16028 16584
rect 14424 16544 15148 16572
rect 15488 16544 16028 16572
rect 14424 16532 14430 16544
rect 14829 16507 14887 16513
rect 14200 16476 14504 16504
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16405 11759 16439
rect 11701 16399 11759 16405
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14476 16445 14504 16476
rect 14829 16473 14841 16507
rect 14875 16504 14887 16507
rect 15488 16504 15516 16544
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16572 17279 16575
rect 17420 16572 17448 16612
rect 17678 16600 17684 16652
rect 17736 16600 17742 16652
rect 18690 16600 18696 16652
rect 18748 16640 18754 16652
rect 19904 16649 19932 16680
rect 20622 16668 20628 16680
rect 20680 16668 20686 16720
rect 20732 16649 20760 16748
rect 22094 16736 22100 16748
rect 22152 16736 22158 16788
rect 19889 16643 19947 16649
rect 18748 16612 19840 16640
rect 18748 16600 18754 16612
rect 17267 16544 17448 16572
rect 17267 16541 17279 16544
rect 17221 16535 17279 16541
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 18782 16572 18788 16584
rect 17644 16544 18788 16572
rect 17644 16532 17650 16544
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 19426 16572 19432 16584
rect 19300 16544 19432 16572
rect 19300 16532 19306 16544
rect 19426 16532 19432 16544
rect 19484 16572 19490 16584
rect 19613 16575 19671 16581
rect 19613 16572 19625 16575
rect 19484 16544 19625 16572
rect 19484 16532 19490 16544
rect 19613 16541 19625 16544
rect 19659 16541 19671 16575
rect 19812 16572 19840 16612
rect 19889 16609 19901 16643
rect 19935 16609 19947 16643
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 19889 16603 19947 16609
rect 19996 16612 20177 16640
rect 19996 16572 20024 16612
rect 20165 16609 20177 16612
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 20717 16643 20775 16649
rect 20717 16609 20729 16643
rect 20763 16609 20775 16643
rect 20717 16603 20775 16609
rect 20990 16600 20996 16652
rect 21048 16600 21054 16652
rect 21542 16600 21548 16652
rect 21600 16640 21606 16652
rect 21600 16612 23428 16640
rect 21600 16600 21606 16612
rect 19812 16544 20024 16572
rect 19613 16535 19671 16541
rect 20346 16532 20352 16584
rect 20404 16532 20410 16584
rect 15562 16513 15568 16516
rect 14875 16476 15516 16504
rect 14875 16473 14887 16476
rect 14829 16467 14887 16473
rect 15556 16467 15568 16513
rect 15562 16464 15568 16467
rect 15620 16464 15626 16516
rect 17034 16504 17040 16516
rect 16684 16476 17040 16504
rect 14369 16439 14427 16445
rect 14369 16436 14381 16439
rect 14332 16408 14381 16436
rect 14332 16396 14338 16408
rect 14369 16405 14381 16408
rect 14415 16405 14427 16439
rect 14369 16399 14427 16405
rect 14461 16439 14519 16445
rect 14461 16405 14473 16439
rect 14507 16405 14519 16439
rect 14461 16399 14519 16405
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 14918 16436 14924 16448
rect 14792 16408 14924 16436
rect 14792 16396 14798 16408
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 16684 16445 16712 16476
rect 17034 16464 17040 16476
rect 17092 16504 17098 16516
rect 17954 16513 17960 16516
rect 17129 16507 17187 16513
rect 17129 16504 17141 16507
rect 17092 16476 17141 16504
rect 17092 16464 17098 16476
rect 17129 16473 17141 16476
rect 17175 16473 17187 16507
rect 17129 16467 17187 16473
rect 17948 16467 17960 16513
rect 17954 16464 17960 16467
rect 18012 16464 18018 16516
rect 20073 16507 20131 16513
rect 20073 16504 20085 16507
rect 18064 16476 20085 16504
rect 16669 16439 16727 16445
rect 16669 16405 16681 16439
rect 16715 16405 16727 16439
rect 16669 16399 16727 16405
rect 16758 16396 16764 16448
rect 16816 16396 16822 16448
rect 17310 16396 17316 16448
rect 17368 16436 17374 16448
rect 18064 16436 18092 16476
rect 20073 16473 20085 16476
rect 20119 16473 20131 16507
rect 20073 16467 20131 16473
rect 21450 16464 21456 16516
rect 21508 16464 21514 16516
rect 23400 16513 23428 16612
rect 22557 16507 22615 16513
rect 22557 16504 22569 16507
rect 22296 16476 22569 16504
rect 17368 16408 18092 16436
rect 17368 16396 17374 16408
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 18414 16436 18420 16448
rect 18196 16408 18420 16436
rect 18196 16396 18202 16408
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 18506 16396 18512 16448
rect 18564 16436 18570 16448
rect 19061 16439 19119 16445
rect 19061 16436 19073 16439
rect 18564 16408 19073 16436
rect 18564 16396 18570 16408
rect 19061 16405 19073 16408
rect 19107 16405 19119 16439
rect 19061 16399 19119 16405
rect 19426 16396 19432 16448
rect 19484 16436 19490 16448
rect 19610 16436 19616 16448
rect 19484 16408 19616 16436
rect 19484 16396 19490 16408
rect 19610 16396 19616 16408
rect 19668 16436 19674 16448
rect 19705 16439 19763 16445
rect 19705 16436 19717 16439
rect 19668 16408 19717 16436
rect 19668 16396 19674 16408
rect 19705 16405 19717 16408
rect 19751 16405 19763 16439
rect 19705 16399 19763 16405
rect 20530 16396 20536 16448
rect 20588 16396 20594 16448
rect 21818 16396 21824 16448
rect 21876 16436 21882 16448
rect 22296 16436 22324 16476
rect 22557 16473 22569 16476
rect 22603 16473 22615 16507
rect 22557 16467 22615 16473
rect 23385 16507 23443 16513
rect 23385 16473 23397 16507
rect 23431 16504 23443 16507
rect 24394 16504 24400 16516
rect 23431 16476 24400 16504
rect 23431 16473 23443 16476
rect 23385 16467 23443 16473
rect 24394 16464 24400 16476
rect 24452 16464 24458 16516
rect 21876 16408 22324 16436
rect 22465 16439 22523 16445
rect 21876 16396 21882 16408
rect 22465 16405 22477 16439
rect 22511 16436 22523 16439
rect 22646 16436 22652 16448
rect 22511 16408 22652 16436
rect 22511 16405 22523 16408
rect 22465 16399 22523 16405
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 1104 16346 26864 16368
rect 1104 16294 3658 16346
rect 3710 16294 3722 16346
rect 3774 16294 3786 16346
rect 3838 16294 3850 16346
rect 3902 16294 3914 16346
rect 3966 16294 3978 16346
rect 4030 16294 7658 16346
rect 7710 16294 7722 16346
rect 7774 16294 7786 16346
rect 7838 16294 7850 16346
rect 7902 16294 7914 16346
rect 7966 16294 7978 16346
rect 8030 16294 11658 16346
rect 11710 16294 11722 16346
rect 11774 16294 11786 16346
rect 11838 16294 11850 16346
rect 11902 16294 11914 16346
rect 11966 16294 11978 16346
rect 12030 16294 15658 16346
rect 15710 16294 15722 16346
rect 15774 16294 15786 16346
rect 15838 16294 15850 16346
rect 15902 16294 15914 16346
rect 15966 16294 15978 16346
rect 16030 16294 19658 16346
rect 19710 16294 19722 16346
rect 19774 16294 19786 16346
rect 19838 16294 19850 16346
rect 19902 16294 19914 16346
rect 19966 16294 19978 16346
rect 20030 16294 23658 16346
rect 23710 16294 23722 16346
rect 23774 16294 23786 16346
rect 23838 16294 23850 16346
rect 23902 16294 23914 16346
rect 23966 16294 23978 16346
rect 24030 16294 26864 16346
rect 1104 16272 26864 16294
rect 2869 16235 2927 16241
rect 2869 16201 2881 16235
rect 2915 16232 2927 16235
rect 3421 16235 3479 16241
rect 2915 16204 3372 16232
rect 2915 16201 2927 16204
rect 2869 16195 2927 16201
rect 2222 16164 2228 16176
rect 1504 16136 2228 16164
rect 1504 16105 1532 16136
rect 2222 16124 2228 16136
rect 2280 16124 2286 16176
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16065 1547 16099
rect 1489 16059 1547 16065
rect 1756 16099 1814 16105
rect 1756 16065 1768 16099
rect 1802 16096 1814 16099
rect 2130 16096 2136 16108
rect 1802 16068 2136 16096
rect 1802 16065 1814 16068
rect 1756 16059 1814 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 3344 16105 3372 16204
rect 3421 16201 3433 16235
rect 3467 16232 3479 16235
rect 4798 16232 4804 16244
rect 3467 16204 4804 16232
rect 3467 16201 3479 16204
rect 3421 16195 3479 16201
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 6638 16192 6644 16244
rect 6696 16192 6702 16244
rect 7098 16192 7104 16244
rect 7156 16232 7162 16244
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 7156 16204 7757 16232
rect 7156 16192 7162 16204
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 7745 16195 7803 16201
rect 7929 16235 7987 16241
rect 7929 16201 7941 16235
rect 7975 16232 7987 16235
rect 8202 16232 8208 16244
rect 7975 16204 8208 16232
rect 7975 16201 7987 16204
rect 7929 16195 7987 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16201 9367 16235
rect 9309 16195 9367 16201
rect 10229 16235 10287 16241
rect 10229 16201 10241 16235
rect 10275 16232 10287 16235
rect 10502 16232 10508 16244
rect 10275 16204 10508 16232
rect 10275 16201 10287 16204
rect 10229 16195 10287 16201
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 5166 16164 5172 16176
rect 4764 16136 5172 16164
rect 4764 16124 4770 16136
rect 5166 16124 5172 16136
rect 5224 16124 5230 16176
rect 5534 16124 5540 16176
rect 5592 16164 5598 16176
rect 6656 16164 6684 16192
rect 5592 16136 6684 16164
rect 5592 16124 5598 16136
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 3375 16068 3740 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 15997 3663 16031
rect 3712 16028 3740 16068
rect 3786 16056 3792 16108
rect 3844 16096 3850 16108
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3844 16068 3985 16096
rect 3844 16056 3850 16068
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 3973 16059 4031 16065
rect 5902 16056 5908 16108
rect 5960 16056 5966 16108
rect 6380 16105 6408 16136
rect 7282 16124 7288 16176
rect 7340 16164 7346 16176
rect 8938 16164 8944 16176
rect 7340 16136 8944 16164
rect 7340 16124 7346 16136
rect 8938 16124 8944 16136
rect 8996 16124 9002 16176
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6621 16099 6679 16105
rect 6621 16096 6633 16099
rect 6365 16059 6423 16065
rect 6472 16068 6633 16096
rect 5166 16028 5172 16040
rect 3712 16000 5172 16028
rect 3605 15991 3663 15997
rect 2774 15920 2780 15972
rect 2832 15960 2838 15972
rect 2961 15963 3019 15969
rect 2961 15960 2973 15963
rect 2832 15932 2973 15960
rect 2832 15920 2838 15932
rect 2961 15929 2973 15932
rect 3007 15929 3019 15963
rect 3620 15960 3648 15991
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 6472 16028 6500 16068
rect 6621 16065 6633 16068
rect 6667 16065 6679 16099
rect 6621 16059 6679 16065
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 7616 16068 8125 16096
rect 7616 16056 7622 16068
rect 8113 16065 8125 16068
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 6104 16000 6500 16028
rect 4154 15960 4160 15972
rect 3620 15932 4160 15960
rect 2961 15923 3019 15929
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 6104 15969 6132 16000
rect 6089 15963 6147 15969
rect 6089 15929 6101 15963
rect 6135 15929 6147 15963
rect 8128 15960 8156 16059
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 8352 16068 8401 16096
rect 8352 16056 8358 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16096 9275 16099
rect 9324 16096 9352 16195
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 10686 16232 10692 16244
rect 10643 16204 10692 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 11072 16204 12434 16232
rect 10042 16124 10048 16176
rect 10100 16164 10106 16176
rect 11072 16164 11100 16204
rect 12406 16164 12434 16204
rect 12618 16192 12624 16244
rect 12676 16232 12682 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 12676 16204 13645 16232
rect 12676 16192 12682 16204
rect 13633 16201 13645 16204
rect 13679 16201 13691 16235
rect 13633 16195 13691 16201
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 14550 16232 14556 16244
rect 14415 16204 14556 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 15562 16192 15568 16244
rect 15620 16232 15626 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15620 16204 15945 16232
rect 15620 16192 15626 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 15933 16195 15991 16201
rect 16758 16192 16764 16244
rect 16816 16192 16822 16244
rect 17310 16192 17316 16244
rect 17368 16192 17374 16244
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 17954 16232 17960 16244
rect 17911 16204 17960 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 18141 16235 18199 16241
rect 18141 16201 18153 16235
rect 18187 16201 18199 16235
rect 18141 16195 18199 16201
rect 10100 16136 11100 16164
rect 11164 16136 12112 16164
rect 12406 16136 13768 16164
rect 10100 16124 10106 16136
rect 9263 16068 9352 16096
rect 9677 16099 9735 16105
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 10318 16096 10324 16108
rect 9723 16068 10324 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 11164 16105 11192 16136
rect 11149 16099 11207 16105
rect 10612 16068 10916 16096
rect 9766 15988 9772 16040
rect 9824 15988 9830 16040
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 16028 10011 16031
rect 10042 16028 10048 16040
rect 9999 16000 10048 16028
rect 9999 15997 10011 16000
rect 9953 15991 10011 15997
rect 10042 15988 10048 16000
rect 10100 16028 10106 16040
rect 10612 16028 10640 16068
rect 10888 16040 10916 16068
rect 11149 16065 11161 16099
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 11422 16056 11428 16108
rect 11480 16096 11486 16108
rect 11957 16099 12015 16105
rect 11957 16096 11969 16099
rect 11480 16068 11969 16096
rect 11480 16056 11486 16068
rect 11957 16065 11969 16068
rect 12003 16065 12015 16099
rect 12084 16096 12112 16136
rect 12084 16068 13216 16096
rect 11957 16059 12015 16065
rect 10100 16000 10640 16028
rect 10689 16031 10747 16037
rect 10100 15988 10106 16000
rect 10689 15997 10701 16031
rect 10735 15997 10747 16031
rect 10689 15991 10747 15997
rect 8128 15932 9628 15960
rect 6089 15923 6147 15929
rect 3326 15852 3332 15904
rect 3384 15892 3390 15904
rect 3789 15895 3847 15901
rect 3789 15892 3801 15895
rect 3384 15864 3801 15892
rect 3384 15852 3390 15864
rect 3789 15861 3801 15864
rect 3835 15861 3847 15895
rect 3789 15855 3847 15861
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 8168 15864 8217 15892
rect 8168 15852 8174 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 9030 15852 9036 15904
rect 9088 15852 9094 15904
rect 9600 15892 9628 15932
rect 10704 15892 10732 15991
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11698 16028 11704 16040
rect 11020 16000 11704 16028
rect 11020 15988 11026 16000
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 11330 15920 11336 15972
rect 11388 15920 11394 15972
rect 12618 15892 12624 15904
rect 9600 15864 12624 15892
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 13078 15852 13084 15904
rect 13136 15852 13142 15904
rect 13188 15901 13216 16068
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 13740 16037 13768 16136
rect 14274 16124 14280 16176
rect 14332 16164 14338 16176
rect 14706 16167 14764 16173
rect 14706 16164 14718 16167
rect 14332 16136 14718 16164
rect 14332 16124 14338 16136
rect 14706 16133 14718 16136
rect 14752 16133 14764 16167
rect 16776 16164 16804 16192
rect 14706 16127 14764 16133
rect 16132 16136 16804 16164
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 15562 16096 15568 16108
rect 14292 16068 15568 16096
rect 13725 16031 13783 16037
rect 13725 15997 13737 16031
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 13998 15988 14004 16040
rect 14056 16028 14062 16040
rect 14292 16028 14320 16068
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 16132 16105 16160 16136
rect 17034 16124 17040 16176
rect 17092 16124 17098 16176
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16065 16175 16099
rect 16117 16059 16175 16065
rect 16666 16056 16672 16108
rect 16724 16056 16730 16108
rect 16850 16105 16856 16108
rect 16817 16099 16856 16105
rect 16817 16065 16829 16099
rect 16817 16059 16856 16065
rect 16850 16056 16856 16059
rect 16908 16056 16914 16108
rect 17218 16105 17224 16108
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17175 16099 17224 16105
rect 17175 16065 17187 16099
rect 17221 16065 17224 16099
rect 17175 16059 17224 16065
rect 14056 16000 14320 16028
rect 14056 15988 14062 16000
rect 14366 15988 14372 16040
rect 14424 16028 14430 16040
rect 14461 16031 14519 16037
rect 14461 16028 14473 16031
rect 14424 16000 14473 16028
rect 14424 15988 14430 16000
rect 14461 15997 14473 16000
rect 14507 15997 14519 16031
rect 16960 16028 16988 16059
rect 17218 16056 17224 16059
rect 17276 16056 17282 16108
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18156 16096 18184 16195
rect 18506 16192 18512 16244
rect 18564 16192 18570 16244
rect 18966 16192 18972 16244
rect 19024 16232 19030 16244
rect 19334 16232 19340 16244
rect 19024 16204 19340 16232
rect 19024 16192 19030 16204
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 19981 16235 20039 16241
rect 19981 16201 19993 16235
rect 20027 16232 20039 16235
rect 20346 16232 20352 16244
rect 20027 16204 20352 16232
rect 20027 16201 20039 16204
rect 19981 16195 20039 16201
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 22830 16192 22836 16244
rect 22888 16232 22894 16244
rect 22925 16235 22983 16241
rect 22925 16232 22937 16235
rect 22888 16204 22937 16232
rect 22888 16192 22894 16204
rect 22925 16201 22937 16204
rect 22971 16201 22983 16235
rect 22925 16195 22983 16201
rect 18782 16164 18788 16176
rect 18095 16068 18184 16096
rect 18708 16136 18788 16164
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 17402 16028 17408 16040
rect 14461 15991 14519 15997
rect 16868 16000 17408 16028
rect 16868 15972 16896 16000
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18414 16028 18420 16040
rect 17920 16000 18420 16028
rect 17920 15988 17926 16000
rect 18414 15988 18420 16000
rect 18472 16028 18478 16040
rect 18708 16037 18736 16136
rect 18782 16124 18788 16136
rect 18840 16124 18846 16176
rect 20530 16164 20536 16176
rect 18984 16136 20536 16164
rect 18984 16105 19012 16136
rect 20530 16124 20536 16136
rect 20588 16124 20594 16176
rect 21818 16124 21824 16176
rect 21876 16124 21882 16176
rect 22554 16124 22560 16176
rect 22612 16124 22618 16176
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16065 19027 16099
rect 18969 16059 19027 16065
rect 19061 16099 19119 16105
rect 19061 16065 19073 16099
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 18601 16031 18659 16037
rect 18601 16028 18613 16031
rect 18472 16000 18613 16028
rect 18472 15988 18478 16000
rect 18601 15997 18613 16000
rect 18647 15997 18659 16031
rect 18601 15991 18659 15997
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 19076 16028 19104 16059
rect 19242 16056 19248 16108
rect 19300 16056 19306 16108
rect 19334 16056 19340 16108
rect 19392 16056 19398 16108
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19576 16068 19625 16096
rect 19576 16056 19582 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16096 19855 16099
rect 20162 16096 20168 16108
rect 19843 16068 20168 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 19812 16028 19840 16059
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 21542 16056 21548 16108
rect 21600 16056 21606 16108
rect 22572 16096 22600 16124
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 22572 16068 23029 16096
rect 23017 16065 23029 16068
rect 23063 16065 23075 16099
rect 23017 16059 23075 16065
rect 26142 16056 26148 16108
rect 26200 16096 26206 16108
rect 26237 16099 26295 16105
rect 26237 16096 26249 16099
rect 26200 16068 26249 16096
rect 26200 16056 26206 16068
rect 26237 16065 26249 16068
rect 26283 16096 26295 16099
rect 26329 16099 26387 16105
rect 26329 16096 26341 16099
rect 26283 16068 26341 16096
rect 26283 16065 26295 16068
rect 26237 16059 26295 16065
rect 26329 16065 26341 16068
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 18840 16000 19104 16028
rect 19168 16000 19840 16028
rect 22066 16000 22569 16028
rect 18840 15988 18846 16000
rect 15841 15963 15899 15969
rect 15841 15929 15853 15963
rect 15887 15960 15899 15963
rect 16114 15960 16120 15972
rect 15887 15932 16120 15960
rect 15887 15929 15899 15932
rect 15841 15923 15899 15929
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 16850 15920 16856 15972
rect 16908 15920 16914 15972
rect 17126 15920 17132 15972
rect 17184 15960 17190 15972
rect 19168 15960 19196 16000
rect 17184 15932 19196 15960
rect 19521 15963 19579 15969
rect 17184 15920 17190 15932
rect 19521 15929 19533 15963
rect 19567 15960 19579 15963
rect 20438 15960 20444 15972
rect 19567 15932 20444 15960
rect 19567 15929 19579 15932
rect 19521 15923 19579 15929
rect 20438 15920 20444 15932
rect 20496 15920 20502 15972
rect 21818 15920 21824 15972
rect 21876 15960 21882 15972
rect 22066 15960 22094 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 21876 15932 22094 15960
rect 21876 15920 21882 15932
rect 13173 15895 13231 15901
rect 13173 15861 13185 15895
rect 13219 15861 13231 15895
rect 13173 15855 13231 15861
rect 14826 15852 14832 15904
rect 14884 15892 14890 15904
rect 18138 15892 18144 15904
rect 14884 15864 18144 15892
rect 14884 15852 14890 15864
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 25958 15852 25964 15904
rect 26016 15892 26022 15904
rect 26145 15895 26203 15901
rect 26145 15892 26157 15895
rect 26016 15864 26157 15892
rect 26016 15852 26022 15864
rect 26145 15861 26157 15864
rect 26191 15861 26203 15895
rect 26145 15855 26203 15861
rect 26234 15852 26240 15904
rect 26292 15892 26298 15904
rect 26421 15895 26479 15901
rect 26421 15892 26433 15895
rect 26292 15864 26433 15892
rect 26292 15852 26298 15864
rect 26421 15861 26433 15864
rect 26467 15861 26479 15895
rect 26421 15855 26479 15861
rect 1104 15802 26864 15824
rect 1104 15750 2918 15802
rect 2970 15750 2982 15802
rect 3034 15750 3046 15802
rect 3098 15750 3110 15802
rect 3162 15750 3174 15802
rect 3226 15750 3238 15802
rect 3290 15750 6918 15802
rect 6970 15750 6982 15802
rect 7034 15750 7046 15802
rect 7098 15750 7110 15802
rect 7162 15750 7174 15802
rect 7226 15750 7238 15802
rect 7290 15750 10918 15802
rect 10970 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 11238 15802
rect 11290 15750 14918 15802
rect 14970 15750 14982 15802
rect 15034 15750 15046 15802
rect 15098 15750 15110 15802
rect 15162 15750 15174 15802
rect 15226 15750 15238 15802
rect 15290 15750 18918 15802
rect 18970 15750 18982 15802
rect 19034 15750 19046 15802
rect 19098 15750 19110 15802
rect 19162 15750 19174 15802
rect 19226 15750 19238 15802
rect 19290 15750 22918 15802
rect 22970 15750 22982 15802
rect 23034 15750 23046 15802
rect 23098 15750 23110 15802
rect 23162 15750 23174 15802
rect 23226 15750 23238 15802
rect 23290 15750 26864 15802
rect 1104 15728 26864 15750
rect 3786 15648 3792 15700
rect 3844 15648 3850 15700
rect 4246 15648 4252 15700
rect 4304 15688 4310 15700
rect 4617 15691 4675 15697
rect 4617 15688 4629 15691
rect 4304 15660 4629 15688
rect 4304 15648 4310 15660
rect 4617 15657 4629 15660
rect 4663 15657 4675 15691
rect 4617 15651 4675 15657
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7374 15688 7380 15700
rect 6972 15660 7380 15688
rect 6972 15648 6978 15660
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 9640 15660 10088 15688
rect 9640 15648 9646 15660
rect 10060 15620 10088 15660
rect 10318 15648 10324 15700
rect 10376 15648 10382 15700
rect 13265 15691 13323 15697
rect 13265 15657 13277 15691
rect 13311 15688 13323 15691
rect 13538 15688 13544 15700
rect 13311 15660 13544 15688
rect 13311 15657 13323 15660
rect 13265 15651 13323 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14829 15691 14887 15697
rect 14829 15688 14841 15691
rect 14240 15660 14841 15688
rect 14240 15648 14246 15660
rect 14829 15657 14841 15660
rect 14875 15657 14887 15691
rect 14829 15651 14887 15657
rect 16114 15648 16120 15700
rect 16172 15688 16178 15700
rect 16482 15688 16488 15700
rect 16172 15660 16488 15688
rect 16172 15648 16178 15660
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 18969 15691 19027 15697
rect 18969 15657 18981 15691
rect 19015 15688 19027 15691
rect 20070 15688 20076 15700
rect 19015 15660 20076 15688
rect 19015 15657 19027 15660
rect 18969 15651 19027 15657
rect 20070 15648 20076 15660
rect 20128 15648 20134 15700
rect 10413 15623 10471 15629
rect 10413 15620 10425 15623
rect 10060 15592 10425 15620
rect 10413 15589 10425 15592
rect 10459 15589 10471 15623
rect 19334 15620 19340 15632
rect 10413 15583 10471 15589
rect 18432 15592 19340 15620
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 5074 15552 5080 15564
rect 4479 15524 5080 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 5534 15512 5540 15564
rect 5592 15512 5598 15564
rect 11698 15512 11704 15564
rect 11756 15552 11762 15564
rect 11885 15555 11943 15561
rect 11885 15552 11897 15555
rect 11756 15524 11897 15552
rect 11756 15512 11762 15524
rect 11885 15521 11897 15524
rect 11931 15521 11943 15555
rect 11885 15515 11943 15521
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15552 15531 15555
rect 15562 15552 15568 15564
rect 15519 15524 15568 15552
rect 15519 15521 15531 15524
rect 15473 15515 15531 15521
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 2222 15444 2228 15496
rect 2280 15444 2286 15496
rect 2492 15487 2550 15493
rect 2492 15453 2504 15487
rect 2538 15484 2550 15487
rect 3326 15484 3332 15496
rect 2538 15456 3332 15484
rect 2538 15453 2550 15456
rect 2492 15447 2550 15453
rect 3326 15444 3332 15456
rect 3384 15444 3390 15496
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4764 15456 4813 15484
rect 4764 15444 4770 15456
rect 4801 15453 4813 15456
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 4982 15444 4988 15496
rect 5040 15444 5046 15496
rect 5166 15444 5172 15496
rect 5224 15444 5230 15496
rect 8110 15444 8116 15496
rect 8168 15493 8174 15496
rect 8168 15484 8180 15493
rect 8389 15487 8447 15493
rect 8168 15456 8213 15484
rect 8168 15447 8180 15456
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8478 15484 8484 15496
rect 8435 15456 8484 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8168 15444 8174 15447
rect 8478 15444 8484 15456
rect 8536 15484 8542 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8536 15456 8953 15484
rect 8536 15444 8542 15456
rect 8941 15453 8953 15456
rect 8987 15484 8999 15487
rect 9674 15484 9680 15496
rect 8987 15456 9680 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10502 15484 10508 15496
rect 9784 15456 10508 15484
rect 4893 15419 4951 15425
rect 4893 15416 4905 15419
rect 4172 15388 4905 15416
rect 4172 15357 4200 15388
rect 4893 15385 4905 15388
rect 4939 15385 4951 15419
rect 4893 15379 4951 15385
rect 5804 15419 5862 15425
rect 5804 15385 5816 15419
rect 5850 15416 5862 15419
rect 5902 15416 5908 15428
rect 5850 15388 5908 15416
rect 5850 15385 5862 15388
rect 5804 15379 5862 15385
rect 5902 15376 5908 15388
rect 5960 15376 5966 15428
rect 7098 15416 7104 15428
rect 6012 15388 7104 15416
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 4157 15351 4215 15357
rect 4157 15348 4169 15351
rect 3651 15320 4169 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 4157 15317 4169 15320
rect 4203 15317 4215 15351
rect 4157 15311 4215 15317
rect 4249 15351 4307 15357
rect 4249 15317 4261 15351
rect 4295 15348 4307 15351
rect 4430 15348 4436 15360
rect 4295 15320 4436 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 4430 15308 4436 15320
rect 4488 15348 4494 15360
rect 6012 15348 6040 15388
rect 7098 15376 7104 15388
rect 7156 15376 7162 15428
rect 9030 15376 9036 15428
rect 9088 15416 9094 15428
rect 9186 15419 9244 15425
rect 9186 15416 9198 15419
rect 9088 15388 9198 15416
rect 9088 15376 9094 15388
rect 9186 15385 9198 15388
rect 9232 15385 9244 15419
rect 9186 15379 9244 15385
rect 4488 15320 6040 15348
rect 4488 15308 4494 15320
rect 7006 15308 7012 15360
rect 7064 15308 7070 15360
rect 8110 15308 8116 15360
rect 8168 15348 8174 15360
rect 9784 15348 9812 15456
rect 10502 15444 10508 15456
rect 10560 15484 10566 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10560 15456 10609 15484
rect 10560 15444 10566 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 10689 15487 10747 15493
rect 10689 15453 10701 15487
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 9858 15376 9864 15428
rect 9916 15416 9922 15428
rect 10704 15416 10732 15447
rect 10870 15444 10876 15496
rect 10928 15444 10934 15496
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 9916 15388 10732 15416
rect 9916 15376 9922 15388
rect 8168 15320 9812 15348
rect 10980 15348 11008 15447
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 12141 15487 12199 15493
rect 12141 15484 12153 15487
rect 11388 15456 12153 15484
rect 11388 15444 11394 15456
rect 12141 15453 12153 15456
rect 12187 15453 12199 15487
rect 14826 15484 14832 15496
rect 12141 15447 12199 15453
rect 12268 15456 14832 15484
rect 12268 15428 12296 15456
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 18432 15493 18460 15592
rect 19334 15580 19340 15592
rect 19392 15580 19398 15632
rect 21174 15620 21180 15632
rect 20732 15592 21180 15620
rect 20732 15561 20760 15592
rect 21174 15580 21180 15592
rect 21232 15620 21238 15632
rect 21542 15620 21548 15632
rect 21232 15592 21548 15620
rect 21232 15580 21238 15592
rect 21542 15580 21548 15592
rect 21600 15580 21606 15632
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15521 20775 15555
rect 20717 15515 20775 15521
rect 24670 15512 24676 15564
rect 24728 15552 24734 15564
rect 26142 15552 26148 15564
rect 24728 15524 26148 15552
rect 24728 15512 24734 15524
rect 26142 15512 26148 15524
rect 26200 15552 26206 15564
rect 26200 15524 26280 15552
rect 26200 15512 26206 15524
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15484 15255 15487
rect 18417 15487 18475 15493
rect 15243 15456 15516 15484
rect 15243 15453 15255 15456
rect 15197 15447 15255 15453
rect 15488 15428 15516 15456
rect 18417 15453 18429 15487
rect 18463 15453 18475 15487
rect 18417 15447 18475 15453
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18564 15456 18705 15484
rect 18564 15444 18570 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 18785 15487 18843 15493
rect 18785 15453 18797 15487
rect 18831 15453 18843 15487
rect 18785 15447 18843 15453
rect 12250 15376 12256 15428
rect 12308 15376 12314 15428
rect 15470 15376 15476 15428
rect 15528 15376 15534 15428
rect 18046 15376 18052 15428
rect 18104 15416 18110 15428
rect 18601 15419 18659 15425
rect 18601 15416 18613 15419
rect 18104 15388 18613 15416
rect 18104 15376 18110 15388
rect 18601 15385 18613 15388
rect 18647 15385 18659 15419
rect 18601 15379 18659 15385
rect 12066 15348 12072 15360
rect 10980 15320 12072 15348
rect 8168 15308 8174 15320
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 14792 15320 15301 15348
rect 14792 15308 14798 15320
rect 15289 15317 15301 15320
rect 15335 15348 15347 15351
rect 17862 15348 17868 15360
rect 15335 15320 17868 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18800 15348 18828 15447
rect 21818 15444 21824 15496
rect 21876 15444 21882 15496
rect 23017 15487 23075 15493
rect 23017 15453 23029 15487
rect 23063 15484 23075 15487
rect 23474 15484 23480 15496
rect 23063 15456 23480 15484
rect 23063 15453 23075 15456
rect 23017 15447 23075 15453
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 24394 15444 24400 15496
rect 24452 15444 24458 15496
rect 26252 15493 26280 15524
rect 26237 15487 26295 15493
rect 26237 15453 26249 15487
rect 26283 15453 26295 15487
rect 26237 15447 26295 15453
rect 20070 15376 20076 15428
rect 20128 15416 20134 15428
rect 20450 15419 20508 15425
rect 20450 15416 20462 15419
rect 20128 15388 20462 15416
rect 20128 15376 20134 15388
rect 20450 15385 20462 15388
rect 20496 15385 20508 15419
rect 20450 15379 20508 15385
rect 24578 15376 24584 15428
rect 24636 15416 24642 15428
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 24636 15388 24685 15416
rect 24636 15376 24642 15388
rect 24673 15385 24685 15388
rect 24719 15385 24731 15419
rect 25958 15416 25964 15428
rect 25898 15388 25964 15416
rect 24673 15379 24731 15385
rect 25958 15376 25964 15388
rect 26016 15376 26022 15428
rect 18012 15320 18828 15348
rect 18012 15308 18018 15320
rect 22830 15308 22836 15360
rect 22888 15348 22894 15360
rect 22925 15351 22983 15357
rect 22925 15348 22937 15351
rect 22888 15320 22937 15348
rect 22888 15308 22894 15320
rect 22925 15317 22937 15320
rect 22971 15317 22983 15351
rect 22925 15311 22983 15317
rect 25038 15308 25044 15360
rect 25096 15348 25102 15360
rect 26145 15351 26203 15357
rect 26145 15348 26157 15351
rect 25096 15320 26157 15348
rect 25096 15308 25102 15320
rect 26145 15317 26157 15320
rect 26191 15317 26203 15351
rect 26145 15311 26203 15317
rect 26326 15308 26332 15360
rect 26384 15308 26390 15360
rect 1104 15258 26864 15280
rect 1104 15206 3658 15258
rect 3710 15206 3722 15258
rect 3774 15206 3786 15258
rect 3838 15206 3850 15258
rect 3902 15206 3914 15258
rect 3966 15206 3978 15258
rect 4030 15206 7658 15258
rect 7710 15206 7722 15258
rect 7774 15206 7786 15258
rect 7838 15206 7850 15258
rect 7902 15206 7914 15258
rect 7966 15206 7978 15258
rect 8030 15206 11658 15258
rect 11710 15206 11722 15258
rect 11774 15206 11786 15258
rect 11838 15206 11850 15258
rect 11902 15206 11914 15258
rect 11966 15206 11978 15258
rect 12030 15206 15658 15258
rect 15710 15206 15722 15258
rect 15774 15206 15786 15258
rect 15838 15206 15850 15258
rect 15902 15206 15914 15258
rect 15966 15206 15978 15258
rect 16030 15206 19658 15258
rect 19710 15206 19722 15258
rect 19774 15206 19786 15258
rect 19838 15206 19850 15258
rect 19902 15206 19914 15258
rect 19966 15206 19978 15258
rect 20030 15206 23658 15258
rect 23710 15206 23722 15258
rect 23774 15206 23786 15258
rect 23838 15206 23850 15258
rect 23902 15206 23914 15258
rect 23966 15206 23978 15258
rect 24030 15206 26864 15258
rect 1104 15184 26864 15206
rect 2130 15104 2136 15156
rect 2188 15104 2194 15156
rect 4249 15147 4307 15153
rect 4249 15113 4261 15147
rect 4295 15144 4307 15147
rect 4338 15144 4344 15156
rect 4295 15116 4344 15144
rect 4295 15113 4307 15116
rect 4249 15107 4307 15113
rect 4338 15104 4344 15116
rect 4396 15144 4402 15156
rect 4709 15147 4767 15153
rect 4709 15144 4721 15147
rect 4396 15116 4721 15144
rect 4396 15104 4402 15116
rect 4709 15113 4721 15116
rect 4755 15113 4767 15147
rect 4709 15107 4767 15113
rect 5902 15104 5908 15156
rect 5960 15104 5966 15156
rect 6733 15147 6791 15153
rect 6733 15113 6745 15147
rect 6779 15144 6791 15147
rect 6914 15144 6920 15156
rect 6779 15116 6920 15144
rect 6779 15113 6791 15116
rect 6733 15107 6791 15113
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 7653 15147 7711 15153
rect 7653 15144 7665 15147
rect 7156 15116 7665 15144
rect 7156 15104 7162 15116
rect 7653 15113 7665 15116
rect 7699 15113 7711 15147
rect 7653 15107 7711 15113
rect 8113 15147 8171 15153
rect 8113 15113 8125 15147
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9858 15104 9864 15156
rect 9916 15104 9922 15156
rect 10318 15144 10324 15156
rect 10244 15116 10324 15144
rect 3136 15079 3194 15085
rect 3136 15045 3148 15079
rect 3182 15076 3194 15079
rect 3326 15076 3332 15088
rect 3182 15048 3332 15076
rect 3182 15045 3194 15048
rect 3136 15039 3194 15045
rect 3326 15036 3332 15048
rect 3384 15036 3390 15088
rect 4154 15036 4160 15088
rect 4212 15076 4218 15088
rect 4212 15048 6868 15076
rect 4212 15036 4218 15048
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 2774 15008 2780 15020
rect 2363 14980 2780 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 2774 14968 2780 14980
rect 2832 14968 2838 15020
rect 6089 15011 6147 15017
rect 6089 14977 6101 15011
rect 6135 15008 6147 15011
rect 6840 15008 6868 15048
rect 8938 15036 8944 15088
rect 8996 15076 9002 15088
rect 10244 15085 10272 15116
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10505 15147 10563 15153
rect 10505 15113 10517 15147
rect 10551 15144 10563 15147
rect 10870 15144 10876 15156
rect 10551 15116 10876 15144
rect 10551 15113 10563 15116
rect 10505 15107 10563 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11422 15144 11428 15156
rect 11112 15116 11428 15144
rect 11112 15104 11118 15116
rect 11422 15104 11428 15116
rect 11480 15144 11486 15156
rect 16850 15144 16856 15156
rect 11480 15116 16856 15144
rect 11480 15104 11486 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 19245 15147 19303 15153
rect 19245 15144 19257 15147
rect 18472 15116 19257 15144
rect 18472 15104 18478 15116
rect 19245 15113 19257 15116
rect 19291 15113 19303 15147
rect 19245 15107 19303 15113
rect 10137 15079 10195 15085
rect 10137 15076 10149 15079
rect 8996 15048 10149 15076
rect 8996 15036 9002 15048
rect 10137 15045 10149 15048
rect 10183 15045 10195 15079
rect 10137 15039 10195 15045
rect 10229 15079 10287 15085
rect 10229 15045 10241 15079
rect 10275 15045 10287 15079
rect 10229 15039 10287 15045
rect 6135 14980 6408 15008
rect 6840 14980 6960 15008
rect 6135 14977 6147 14980
rect 6089 14971 6147 14977
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2869 14943 2927 14949
rect 2869 14940 2881 14943
rect 2280 14912 2881 14940
rect 2280 14900 2286 14912
rect 2869 14909 2881 14912
rect 2915 14909 2927 14943
rect 2869 14903 2927 14909
rect 4798 14900 4804 14952
rect 4856 14900 4862 14952
rect 4890 14900 4896 14952
rect 4948 14900 4954 14952
rect 4338 14764 4344 14816
rect 4396 14764 4402 14816
rect 4816 14804 4844 14900
rect 6380 14881 6408 14980
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 6932 14949 6960 14980
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7742 15008 7748 15020
rect 7064 14980 7748 15008
rect 7064 14968 7070 14980
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 8202 14968 8208 15020
rect 8260 14968 8266 15020
rect 8478 14968 8484 15020
rect 8536 15017 8542 15020
rect 8754 15017 8760 15020
rect 8536 15008 8546 15017
rect 8748 15008 8760 15017
rect 8536 14980 8581 15008
rect 8715 14980 8760 15008
rect 8536 14971 8546 14980
rect 8748 14971 8760 14980
rect 8536 14968 8542 14971
rect 8754 14968 8760 14971
rect 8812 14968 8818 15020
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 9088 14980 9965 15008
rect 9088 14968 9094 14980
rect 9953 14977 9965 14980
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 7466 14900 7472 14952
rect 7524 14900 7530 14952
rect 6365 14875 6423 14881
rect 6365 14841 6377 14875
rect 6411 14841 6423 14875
rect 6840 14872 6868 14900
rect 7558 14872 7564 14884
rect 6840 14844 7564 14872
rect 6365 14835 6423 14841
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 8389 14875 8447 14881
rect 8389 14841 8401 14875
rect 8435 14872 8447 14875
rect 8478 14872 8484 14884
rect 8435 14844 8484 14872
rect 8435 14841 8447 14844
rect 8389 14835 8447 14841
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 10152 14872 10180 15039
rect 13998 15036 14004 15088
rect 14056 15036 14062 15088
rect 17862 15036 17868 15088
rect 17920 15076 17926 15088
rect 18598 15076 18604 15088
rect 17920 15048 18604 15076
rect 17920 15036 17926 15048
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 10594 15008 10600 15020
rect 10367 14980 10600 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 19260 15008 19288 15107
rect 19334 15104 19340 15156
rect 19392 15104 19398 15156
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15113 19763 15147
rect 19705 15107 19763 15113
rect 19981 15147 20039 15153
rect 19981 15113 19993 15147
rect 20027 15144 20039 15147
rect 20070 15144 20076 15156
rect 20027 15116 20076 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 19334 15008 19340 15020
rect 19260 14980 19340 15008
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19720 15008 19748 15107
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 22830 15036 22836 15088
rect 22888 15036 22894 15088
rect 19797 15011 19855 15017
rect 19797 15008 19809 15011
rect 19720 14980 19809 15008
rect 19797 14977 19809 14980
rect 19843 14977 19855 15011
rect 19797 14971 19855 14977
rect 24118 14968 24124 15020
rect 24176 15008 24182 15020
rect 24670 15008 24676 15020
rect 24176 14980 24676 15008
rect 24176 14968 24182 14980
rect 24670 14968 24676 14980
rect 24728 15008 24734 15020
rect 25041 15011 25099 15017
rect 25041 15008 25053 15011
rect 24728 14980 25053 15008
rect 24728 14968 24734 14980
rect 25041 14977 25053 14980
rect 25087 14977 25099 15011
rect 25041 14971 25099 14977
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14909 19211 14943
rect 19153 14903 19211 14909
rect 17678 14872 17684 14884
rect 10152 14844 17684 14872
rect 17678 14832 17684 14844
rect 17736 14832 17742 14884
rect 19168 14872 19196 14903
rect 21818 14900 21824 14952
rect 21876 14900 21882 14952
rect 22097 14943 22155 14949
rect 22097 14909 22109 14943
rect 22143 14940 22155 14943
rect 24210 14940 24216 14952
rect 22143 14912 24216 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 24210 14900 24216 14912
rect 24268 14900 24274 14952
rect 25593 14943 25651 14949
rect 25593 14909 25605 14943
rect 25639 14940 25651 14943
rect 25958 14940 25964 14952
rect 25639 14912 25964 14940
rect 25639 14909 25651 14912
rect 25593 14903 25651 14909
rect 25958 14900 25964 14912
rect 26016 14900 26022 14952
rect 20438 14872 20444 14884
rect 19168 14844 20444 14872
rect 20438 14832 20444 14844
rect 20496 14832 20502 14884
rect 9766 14804 9772 14816
rect 4816 14776 9772 14804
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 15289 14807 15347 14813
rect 15289 14804 15301 14807
rect 14884 14776 15301 14804
rect 14884 14764 14890 14776
rect 15289 14773 15301 14776
rect 15335 14773 15347 14807
rect 15289 14767 15347 14773
rect 23569 14807 23627 14813
rect 23569 14773 23581 14807
rect 23615 14804 23627 14807
rect 24670 14804 24676 14816
rect 23615 14776 24676 14804
rect 23615 14773 23627 14776
rect 23569 14767 23627 14773
rect 24670 14764 24676 14776
rect 24728 14764 24734 14816
rect 25130 14764 25136 14816
rect 25188 14764 25194 14816
rect 26418 14764 26424 14816
rect 26476 14804 26482 14816
rect 26513 14807 26571 14813
rect 26513 14804 26525 14807
rect 26476 14776 26525 14804
rect 26476 14764 26482 14776
rect 26513 14773 26525 14776
rect 26559 14773 26571 14807
rect 26513 14767 26571 14773
rect 1104 14714 26864 14736
rect 1104 14662 2918 14714
rect 2970 14662 2982 14714
rect 3034 14662 3046 14714
rect 3098 14662 3110 14714
rect 3162 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 6918 14714
rect 6970 14662 6982 14714
rect 7034 14662 7046 14714
rect 7098 14662 7110 14714
rect 7162 14662 7174 14714
rect 7226 14662 7238 14714
rect 7290 14662 10918 14714
rect 10970 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 11238 14714
rect 11290 14662 14918 14714
rect 14970 14662 14982 14714
rect 15034 14662 15046 14714
rect 15098 14662 15110 14714
rect 15162 14662 15174 14714
rect 15226 14662 15238 14714
rect 15290 14662 18918 14714
rect 18970 14662 18982 14714
rect 19034 14662 19046 14714
rect 19098 14662 19110 14714
rect 19162 14662 19174 14714
rect 19226 14662 19238 14714
rect 19290 14662 22918 14714
rect 22970 14662 22982 14714
rect 23034 14662 23046 14714
rect 23098 14662 23110 14714
rect 23162 14662 23174 14714
rect 23226 14662 23238 14714
rect 23290 14662 26864 14714
rect 1104 14640 26864 14662
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 3326 14600 3332 14612
rect 3283 14572 3332 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 6270 14560 6276 14612
rect 6328 14600 6334 14612
rect 6822 14600 6828 14612
rect 6328 14572 6828 14600
rect 6328 14560 6334 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 8260 14572 9045 14600
rect 8260 14560 8266 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9033 14563 9091 14569
rect 13722 14560 13728 14612
rect 13780 14560 13786 14612
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 18782 14600 18788 14612
rect 16807 14572 18788 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19334 14560 19340 14612
rect 19392 14560 19398 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 26329 14603 26387 14609
rect 26329 14600 26341 14603
rect 19484 14572 26341 14600
rect 19484 14560 19490 14572
rect 6730 14492 6736 14544
rect 6788 14532 6794 14544
rect 7466 14532 7472 14544
rect 6788 14504 7472 14532
rect 6788 14492 6794 14504
rect 7466 14492 7472 14504
rect 7524 14532 7530 14544
rect 7524 14504 12020 14532
rect 7524 14492 7530 14504
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 11992 14464 12020 14504
rect 12066 14492 12072 14544
rect 12124 14532 12130 14544
rect 13740 14532 13768 14560
rect 18325 14535 18383 14541
rect 12124 14504 16252 14532
rect 12124 14492 12130 14504
rect 12710 14464 12716 14476
rect 11992 14436 12716 14464
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13722 14464 13728 14476
rect 13504 14436 13728 14464
rect 13504 14424 13510 14436
rect 13722 14424 13728 14436
rect 13780 14464 13786 14476
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 13780 14436 15117 14464
rect 13780 14424 13786 14436
rect 15105 14433 15117 14436
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 4338 14396 4344 14408
rect 3467 14368 4344 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14396 9459 14399
rect 9858 14396 9864 14408
rect 9447 14368 9864 14396
rect 9447 14365 9459 14368
rect 9401 14359 9459 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 14507 14368 14596 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 9766 14328 9772 14340
rect 9539 14300 9772 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 14274 14220 14280 14272
rect 14332 14220 14338 14272
rect 14568 14269 14596 14368
rect 15378 14356 15384 14408
rect 15436 14356 15442 14408
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 15488 14368 15669 14396
rect 14921 14331 14979 14337
rect 14921 14297 14933 14331
rect 14967 14328 14979 14331
rect 15102 14328 15108 14340
rect 14967 14300 15108 14328
rect 14967 14297 14979 14300
rect 14921 14291 14979 14297
rect 15102 14288 15108 14300
rect 15160 14328 15166 14340
rect 15488 14328 15516 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 15746 14356 15752 14408
rect 15804 14356 15810 14408
rect 16224 14405 16252 14504
rect 18325 14501 18337 14535
rect 18371 14532 18383 14535
rect 18690 14532 18696 14544
rect 18371 14504 18696 14532
rect 18371 14501 18383 14504
rect 18325 14495 18383 14501
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14365 16359 14399
rect 16301 14359 16359 14365
rect 15160 14300 15516 14328
rect 15565 14331 15623 14337
rect 15160 14288 15166 14300
rect 15565 14297 15577 14331
rect 15611 14297 15623 14331
rect 16316 14328 16344 14359
rect 16482 14356 16488 14408
rect 16540 14356 16546 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 16666 14396 16672 14408
rect 16623 14368 16672 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 16666 14356 16672 14368
rect 16724 14396 16730 14408
rect 16942 14396 16948 14408
rect 16724 14368 16948 14396
rect 16724 14356 16730 14368
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 18463 14399 18521 14405
rect 18463 14396 18475 14399
rect 17644 14368 18475 14396
rect 17644 14356 17650 14368
rect 18463 14365 18475 14368
rect 18509 14365 18521 14399
rect 18463 14359 18521 14365
rect 18690 14356 18696 14408
rect 18748 14356 18754 14408
rect 18874 14396 18880 14408
rect 18835 14368 18880 14396
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 19536 14405 19564 14572
rect 26329 14569 26341 14572
rect 26375 14569 26387 14603
rect 26329 14563 26387 14569
rect 21174 14424 21180 14476
rect 21232 14424 21238 14476
rect 21453 14467 21511 14473
rect 21453 14433 21465 14467
rect 21499 14464 21511 14467
rect 23566 14464 23572 14476
rect 21499 14436 23572 14464
rect 21499 14433 21511 14436
rect 21453 14427 21511 14433
rect 23566 14424 23572 14436
rect 23624 14424 23630 14476
rect 24670 14424 24676 14476
rect 24728 14424 24734 14476
rect 18969 14399 19027 14405
rect 18969 14365 18981 14399
rect 19015 14365 19027 14399
rect 18969 14359 19027 14365
rect 19521 14399 19579 14405
rect 19521 14365 19533 14399
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 23474 14396 23480 14408
rect 23247 14368 23480 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 15565 14291 15623 14297
rect 15948 14300 16344 14328
rect 14553 14263 14611 14269
rect 14553 14229 14565 14263
rect 14599 14229 14611 14263
rect 14553 14223 14611 14229
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14884 14232 15025 14260
rect 14884 14220 14890 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 15470 14220 15476 14272
rect 15528 14260 15534 14272
rect 15580 14260 15608 14291
rect 15948 14269 15976 14300
rect 18598 14288 18604 14340
rect 18656 14288 18662 14340
rect 15528 14232 15608 14260
rect 15933 14263 15991 14269
rect 15528 14220 15534 14232
rect 15933 14229 15945 14263
rect 15979 14229 15991 14263
rect 15933 14223 15991 14229
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 18984 14260 19012 14359
rect 23474 14356 23480 14368
rect 23532 14396 23538 14408
rect 24118 14396 24124 14408
rect 23532 14368 24124 14396
rect 23532 14356 23538 14368
rect 24118 14356 24124 14368
rect 24176 14356 24182 14408
rect 24394 14356 24400 14408
rect 24452 14356 24458 14408
rect 26418 14356 26424 14408
rect 26476 14356 26482 14408
rect 23109 14331 23167 14337
rect 23109 14328 23121 14331
rect 22678 14300 23121 14328
rect 23109 14297 23121 14300
rect 23155 14297 23167 14331
rect 23109 14291 23167 14297
rect 25130 14288 25136 14340
rect 25188 14288 25194 14340
rect 18840 14232 19012 14260
rect 18840 14220 18846 14232
rect 22278 14220 22284 14272
rect 22336 14260 22342 14272
rect 22925 14263 22983 14269
rect 22925 14260 22937 14263
rect 22336 14232 22937 14260
rect 22336 14220 22342 14232
rect 22925 14229 22937 14232
rect 22971 14229 22983 14263
rect 22925 14223 22983 14229
rect 24854 14220 24860 14272
rect 24912 14260 24918 14272
rect 26145 14263 26203 14269
rect 26145 14260 26157 14263
rect 24912 14232 26157 14260
rect 24912 14220 24918 14232
rect 26145 14229 26157 14232
rect 26191 14229 26203 14263
rect 26145 14223 26203 14229
rect 1104 14170 26864 14192
rect 1104 14118 3658 14170
rect 3710 14118 3722 14170
rect 3774 14118 3786 14170
rect 3838 14118 3850 14170
rect 3902 14118 3914 14170
rect 3966 14118 3978 14170
rect 4030 14118 7658 14170
rect 7710 14118 7722 14170
rect 7774 14118 7786 14170
rect 7838 14118 7850 14170
rect 7902 14118 7914 14170
rect 7966 14118 7978 14170
rect 8030 14118 11658 14170
rect 11710 14118 11722 14170
rect 11774 14118 11786 14170
rect 11838 14118 11850 14170
rect 11902 14118 11914 14170
rect 11966 14118 11978 14170
rect 12030 14118 15658 14170
rect 15710 14118 15722 14170
rect 15774 14118 15786 14170
rect 15838 14118 15850 14170
rect 15902 14118 15914 14170
rect 15966 14118 15978 14170
rect 16030 14118 19658 14170
rect 19710 14118 19722 14170
rect 19774 14118 19786 14170
rect 19838 14118 19850 14170
rect 19902 14118 19914 14170
rect 19966 14118 19978 14170
rect 20030 14118 23658 14170
rect 23710 14118 23722 14170
rect 23774 14118 23786 14170
rect 23838 14118 23850 14170
rect 23902 14118 23914 14170
rect 23966 14118 23978 14170
rect 24030 14118 26864 14170
rect 1104 14096 26864 14118
rect 13541 14059 13599 14065
rect 9646 14028 11100 14056
rect 7374 13948 7380 14000
rect 7432 13988 7438 14000
rect 9646 13988 9674 14028
rect 7432 13960 9674 13988
rect 7432 13948 7438 13960
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 10612 13852 10640 13883
rect 10686 13880 10692 13932
rect 10744 13880 10750 13932
rect 10873 13923 10931 13929
rect 10873 13889 10885 13923
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 10975 13923 11033 13929
rect 10975 13889 10987 13923
rect 11021 13920 11033 13923
rect 11072 13920 11100 14028
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 14182 14056 14188 14068
rect 13587 14028 14188 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 15013 14059 15071 14065
rect 15013 14025 15025 14059
rect 15059 14056 15071 14059
rect 15102 14056 15108 14068
rect 15059 14028 15108 14056
rect 15059 14025 15071 14028
rect 15013 14019 15071 14025
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 17037 14059 17095 14065
rect 17037 14056 17049 14059
rect 16540 14028 17049 14056
rect 16540 14016 16546 14028
rect 17037 14025 17049 14028
rect 17083 14025 17095 14059
rect 17037 14019 17095 14025
rect 18785 14059 18843 14065
rect 18785 14025 18797 14059
rect 18831 14056 18843 14059
rect 18874 14056 18880 14068
rect 18831 14028 18880 14056
rect 18831 14025 18843 14028
rect 18785 14019 18843 14025
rect 18874 14016 18880 14028
rect 18932 14056 18938 14068
rect 19245 14059 19303 14065
rect 19245 14056 19257 14059
rect 18932 14028 19257 14056
rect 18932 14016 18938 14028
rect 19245 14025 19257 14028
rect 19291 14025 19303 14059
rect 19245 14019 19303 14025
rect 13900 13991 13958 13997
rect 13900 13957 13912 13991
rect 13946 13988 13958 13991
rect 14274 13988 14280 14000
rect 13946 13960 14280 13988
rect 13946 13957 13958 13960
rect 13900 13951 13958 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 17865 13991 17923 13997
rect 17865 13957 17877 13991
rect 17911 13988 17923 13991
rect 18046 13988 18052 14000
rect 17911 13960 18052 13988
rect 17911 13957 17923 13960
rect 17865 13951 17923 13957
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 18690 13948 18696 14000
rect 18748 13948 18754 14000
rect 22278 13948 22284 14000
rect 22336 13948 22342 14000
rect 22830 13948 22836 14000
rect 22888 13948 22894 14000
rect 24213 13991 24271 13997
rect 24213 13957 24225 13991
rect 24259 13988 24271 13991
rect 24946 13988 24952 14000
rect 24259 13960 24952 13988
rect 24259 13957 24271 13960
rect 24213 13951 24271 13957
rect 24946 13948 24952 13960
rect 25004 13948 25010 14000
rect 26326 13988 26332 14000
rect 25898 13960 26332 13988
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 11021 13892 11100 13920
rect 11021 13889 11033 13892
rect 10975 13883 11033 13889
rect 10888 13882 10928 13883
rect 10900 13852 10928 13882
rect 11422 13880 11428 13932
rect 11480 13920 11486 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11480 13892 11713 13920
rect 11480 13880 11486 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11790 13880 11796 13932
rect 11848 13880 11854 13932
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 9824 13824 10732 13852
rect 10900 13824 11529 13852
rect 9824 13812 9830 13824
rect 10410 13744 10416 13796
rect 10468 13744 10474 13796
rect 10704 13784 10732 13824
rect 11517 13821 11529 13824
rect 11563 13821 11575 13855
rect 11992 13852 12020 13883
rect 12066 13880 12072 13932
rect 12124 13880 12130 13932
rect 12158 13880 12164 13932
rect 12216 13880 12222 13932
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 14458 13920 14464 13932
rect 13403 13892 14464 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 15372 13923 15430 13929
rect 15372 13889 15384 13923
rect 15418 13920 15430 13923
rect 15746 13920 15752 13932
rect 15418 13892 15752 13920
rect 15418 13889 15430 13892
rect 15372 13883 15430 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 17175 13892 17969 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17957 13889 17969 13892
rect 18003 13920 18015 13923
rect 18708 13920 18736 13948
rect 19426 13920 19432 13932
rect 18003 13892 19432 13920
rect 18003 13889 18015 13892
rect 17957 13883 18015 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 20070 13880 20076 13932
rect 20128 13920 20134 13932
rect 20358 13923 20416 13929
rect 20358 13920 20370 13923
rect 20128 13892 20370 13920
rect 20128 13880 20134 13892
rect 20358 13889 20370 13892
rect 20404 13889 20416 13923
rect 20358 13883 20416 13889
rect 24118 13880 24124 13932
rect 24176 13880 24182 13932
rect 12250 13852 12256 13864
rect 11992 13824 12256 13852
rect 11517 13815 11575 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13821 13691 13855
rect 13633 13815 13691 13821
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13821 15163 13855
rect 15105 13815 15163 13821
rect 17221 13855 17279 13861
rect 17221 13821 17233 13855
rect 17267 13821 17279 13855
rect 17221 13815 17279 13821
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18509 13855 18567 13861
rect 18509 13821 18521 13855
rect 18555 13821 18567 13855
rect 18509 13815 18567 13821
rect 18693 13855 18751 13861
rect 18693 13821 18705 13855
rect 18739 13852 18751 13855
rect 19334 13852 19340 13864
rect 18739 13824 19340 13852
rect 18739 13821 18751 13824
rect 18693 13815 18751 13821
rect 13538 13784 13544 13796
rect 10704 13756 13544 13784
rect 13538 13744 13544 13756
rect 13596 13744 13602 13796
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 5258 13716 5264 13728
rect 4856 13688 5264 13716
rect 4856 13676 4862 13688
rect 5258 13676 5264 13688
rect 5316 13716 5322 13728
rect 11330 13716 11336 13728
rect 5316 13688 11336 13716
rect 5316 13676 5322 13688
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 12345 13719 12403 13725
rect 12345 13685 12357 13719
rect 12391 13716 12403 13719
rect 12526 13716 12532 13728
rect 12391 13688 12532 13716
rect 12391 13685 12403 13688
rect 12345 13679 12403 13685
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 13648 13716 13676 13815
rect 13814 13716 13820 13728
rect 13648 13688 13820 13716
rect 13814 13676 13820 13688
rect 13872 13716 13878 13728
rect 14366 13716 14372 13728
rect 13872 13688 14372 13716
rect 13872 13676 13878 13688
rect 14366 13676 14372 13688
rect 14424 13716 14430 13728
rect 15120 13716 15148 13815
rect 16850 13744 16856 13796
rect 16908 13784 16914 13796
rect 17236 13784 17264 13815
rect 16908 13756 17264 13784
rect 16908 13744 16914 13756
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 18064 13784 18092 13815
rect 17368 13756 18092 13784
rect 17368 13744 17374 13756
rect 18414 13744 18420 13796
rect 18472 13784 18478 13796
rect 18524 13784 18552 13815
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13852 20683 13855
rect 20714 13852 20720 13864
rect 20671 13824 20720 13852
rect 20671 13821 20683 13824
rect 20625 13815 20683 13821
rect 20714 13812 20720 13824
rect 20772 13852 20778 13864
rect 21818 13852 21824 13864
rect 20772 13824 21824 13852
rect 20772 13812 20778 13824
rect 21818 13812 21824 13824
rect 21876 13852 21882 13864
rect 22002 13852 22008 13864
rect 21876 13824 22008 13852
rect 21876 13812 21882 13824
rect 22002 13812 22008 13824
rect 22060 13812 22066 13864
rect 23474 13812 23480 13864
rect 23532 13852 23538 13864
rect 23753 13855 23811 13861
rect 23753 13852 23765 13855
rect 23532 13824 23765 13852
rect 23532 13812 23538 13824
rect 23753 13821 23765 13824
rect 23799 13821 23811 13855
rect 23753 13815 23811 13821
rect 24394 13812 24400 13864
rect 24452 13812 24458 13864
rect 18472 13756 18552 13784
rect 18472 13744 18478 13756
rect 14424 13688 15148 13716
rect 14424 13676 14430 13688
rect 15838 13676 15844 13728
rect 15896 13716 15902 13728
rect 16669 13719 16727 13725
rect 16669 13716 16681 13719
rect 15896 13688 16681 13716
rect 15896 13676 15902 13688
rect 16669 13685 16681 13688
rect 16715 13685 16727 13719
rect 16669 13679 16727 13685
rect 16942 13676 16948 13728
rect 17000 13716 17006 13728
rect 17497 13719 17555 13725
rect 17497 13716 17509 13719
rect 17000 13688 17509 13716
rect 17000 13676 17006 13688
rect 17497 13685 17509 13688
rect 17543 13685 17555 13719
rect 17497 13679 17555 13685
rect 19153 13719 19211 13725
rect 19153 13685 19165 13719
rect 19199 13716 19211 13719
rect 19518 13716 19524 13728
rect 19199 13688 19524 13716
rect 19199 13685 19211 13688
rect 19153 13679 19211 13685
rect 19518 13676 19524 13688
rect 19576 13676 19582 13728
rect 24660 13719 24718 13725
rect 24660 13685 24672 13719
rect 24706 13716 24718 13719
rect 25222 13716 25228 13728
rect 24706 13688 25228 13716
rect 24706 13685 24718 13688
rect 24660 13679 24718 13685
rect 25222 13676 25228 13688
rect 25280 13676 25286 13728
rect 26142 13676 26148 13728
rect 26200 13676 26206 13728
rect 1104 13626 26864 13648
rect 1104 13574 2918 13626
rect 2970 13574 2982 13626
rect 3034 13574 3046 13626
rect 3098 13574 3110 13626
rect 3162 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 6918 13626
rect 6970 13574 6982 13626
rect 7034 13574 7046 13626
rect 7098 13574 7110 13626
rect 7162 13574 7174 13626
rect 7226 13574 7238 13626
rect 7290 13574 10918 13626
rect 10970 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 11238 13626
rect 11290 13574 14918 13626
rect 14970 13574 14982 13626
rect 15034 13574 15046 13626
rect 15098 13574 15110 13626
rect 15162 13574 15174 13626
rect 15226 13574 15238 13626
rect 15290 13574 18918 13626
rect 18970 13574 18982 13626
rect 19034 13574 19046 13626
rect 19098 13574 19110 13626
rect 19162 13574 19174 13626
rect 19226 13574 19238 13626
rect 19290 13574 22918 13626
rect 22970 13574 22982 13626
rect 23034 13574 23046 13626
rect 23098 13574 23110 13626
rect 23162 13574 23174 13626
rect 23226 13574 23238 13626
rect 23290 13574 26864 13626
rect 1104 13552 26864 13574
rect 5905 13515 5963 13521
rect 4356 13484 5856 13512
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 4062 13376 4068 13388
rect 1995 13348 4068 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 4062 13336 4068 13348
rect 4120 13376 4126 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4120 13348 4261 13376
rect 4120 13336 4126 13348
rect 4249 13345 4261 13348
rect 4295 13376 4307 13379
rect 4356 13376 4384 13484
rect 4890 13444 4896 13456
rect 4448 13416 4896 13444
rect 4448 13388 4476 13416
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 5261 13447 5319 13453
rect 5261 13413 5273 13447
rect 5307 13444 5319 13447
rect 5307 13416 5764 13444
rect 5307 13413 5319 13416
rect 5261 13407 5319 13413
rect 4295 13348 4384 13376
rect 4295 13345 4307 13348
rect 4249 13339 4307 13345
rect 4430 13336 4436 13388
rect 4488 13336 4494 13388
rect 4982 13336 4988 13388
rect 5040 13336 5046 13388
rect 5736 13385 5764 13416
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13345 5779 13379
rect 5828 13376 5856 13484
rect 5905 13481 5917 13515
rect 5951 13512 5963 13515
rect 7558 13512 7564 13524
rect 5951 13484 7564 13512
rect 5951 13481 5963 13484
rect 5905 13475 5963 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 11425 13515 11483 13521
rect 11425 13481 11437 13515
rect 11471 13512 11483 13515
rect 11514 13512 11520 13524
rect 11471 13484 11520 13512
rect 11471 13481 11483 13484
rect 11425 13475 11483 13481
rect 11514 13472 11520 13484
rect 11572 13512 11578 13524
rect 11790 13512 11796 13524
rect 11572 13484 11796 13512
rect 11572 13472 11578 13484
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 15436 13484 15485 13512
rect 15436 13472 15442 13484
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 15473 13475 15531 13481
rect 15746 13472 15752 13524
rect 15804 13472 15810 13524
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 18414 13512 18420 13524
rect 16264 13484 18420 13512
rect 16264 13472 16270 13484
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 18782 13472 18788 13524
rect 18840 13512 18846 13524
rect 19061 13515 19119 13521
rect 19061 13512 19073 13515
rect 18840 13484 19073 13512
rect 18840 13472 18846 13484
rect 19061 13481 19073 13484
rect 19107 13481 19119 13515
rect 19061 13475 19119 13481
rect 22830 13472 22836 13524
rect 22888 13512 22894 13524
rect 23017 13515 23075 13521
rect 23017 13512 23029 13515
rect 22888 13484 23029 13512
rect 22888 13472 22894 13484
rect 23017 13481 23029 13484
rect 23063 13481 23075 13515
rect 23017 13475 23075 13481
rect 6089 13447 6147 13453
rect 6089 13413 6101 13447
rect 6135 13444 6147 13447
rect 7374 13444 7380 13456
rect 6135 13416 7380 13444
rect 6135 13413 6147 13416
rect 6089 13407 6147 13413
rect 7374 13404 7380 13416
rect 7432 13404 7438 13456
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 8938 13444 8944 13456
rect 8352 13416 8944 13444
rect 8352 13404 8358 13416
rect 8938 13404 8944 13416
rect 8996 13404 9002 13456
rect 9490 13404 9496 13456
rect 9548 13444 9554 13456
rect 10873 13447 10931 13453
rect 9548 13416 9720 13444
rect 9548 13404 9554 13416
rect 5828 13348 7052 13376
rect 5721 13339 5779 13345
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 2096 13280 2237 13308
rect 2096 13268 2102 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 2700 13240 2728 13271
rect 2958 13268 2964 13320
rect 3016 13268 3022 13320
rect 4522 13268 4528 13320
rect 4580 13308 4586 13320
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4580 13280 4629 13308
rect 4580 13268 4586 13280
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 4710 13311 4768 13317
rect 4710 13277 4722 13311
rect 4756 13277 4768 13311
rect 4710 13271 4768 13277
rect 4724 13240 4752 13271
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4856 13280 4905 13308
rect 4856 13268 4862 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 5000 13308 5028 13336
rect 5082 13311 5140 13317
rect 5082 13308 5094 13311
rect 5000 13280 5094 13308
rect 4893 13271 4951 13277
rect 5082 13277 5094 13280
rect 5128 13277 5140 13311
rect 5082 13271 5140 13277
rect 5626 13268 5632 13320
rect 5684 13268 5690 13320
rect 5902 13268 5908 13320
rect 5960 13268 5966 13320
rect 6178 13268 6184 13320
rect 6236 13268 6242 13320
rect 7024 13249 7052 13348
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7193 13379 7251 13385
rect 7193 13376 7205 13379
rect 7156 13348 7205 13376
rect 7156 13336 7162 13348
rect 7193 13345 7205 13348
rect 7239 13376 7251 13379
rect 9582 13376 9588 13388
rect 7239 13348 9588 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 9582 13336 9588 13348
rect 9640 13336 9646 13388
rect 9692 13385 9720 13416
rect 10873 13413 10885 13447
rect 10919 13413 10931 13447
rect 10873 13407 10931 13413
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10008 13348 10241 13376
rect 10008 13336 10014 13348
rect 10229 13345 10241 13348
rect 10275 13376 10287 13379
rect 10594 13376 10600 13388
rect 10275 13348 10600 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 10686 13308 10692 13320
rect 10551 13280 10692 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 10888 13308 10916 13407
rect 18598 13404 18604 13456
rect 18656 13444 18662 13456
rect 19242 13444 19248 13456
rect 18656 13416 19248 13444
rect 18656 13404 18662 13416
rect 19242 13404 19248 13416
rect 19300 13404 19306 13456
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13376 12863 13379
rect 13814 13376 13820 13388
rect 12851 13348 13820 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 13814 13336 13820 13348
rect 13872 13376 13878 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13872 13348 14105 13376
rect 13872 13336 13878 13348
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 14093 13339 14151 13345
rect 15396 13348 17049 13376
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10888 13280 10977 13308
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 12526 13268 12532 13320
rect 12584 13317 12590 13320
rect 12584 13271 12596 13317
rect 12584 13268 12590 13271
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 14108 13308 14136 13339
rect 15396 13308 15424 13348
rect 17037 13345 17049 13348
rect 17083 13345 17095 13379
rect 17037 13339 17095 13345
rect 18230 13336 18236 13388
rect 18288 13376 18294 13388
rect 18288 13348 18920 13376
rect 18288 13336 18294 13348
rect 14108 13280 15424 13308
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15896 13280 15945 13308
rect 15896 13268 15902 13280
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 16482 13268 16488 13320
rect 16540 13268 16546 13320
rect 16666 13308 16672 13320
rect 16592 13280 16672 13308
rect 4985 13243 5043 13249
rect 4985 13240 4997 13243
rect 2700 13212 3832 13240
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 2188 13144 2513 13172
rect 2188 13132 2194 13144
rect 2501 13141 2513 13144
rect 2547 13141 2559 13175
rect 2501 13135 2559 13141
rect 2774 13132 2780 13184
rect 2832 13132 2838 13184
rect 3804 13181 3832 13212
rect 4172 13212 4752 13240
rect 4816 13212 4997 13240
rect 4172 13184 4200 13212
rect 4816 13184 4844 13212
rect 4985 13209 4997 13212
rect 5031 13209 5043 13243
rect 4985 13203 5043 13209
rect 7009 13243 7067 13249
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 9493 13243 9551 13249
rect 7055 13212 9260 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 3789 13175 3847 13181
rect 3789 13141 3801 13175
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 4154 13132 4160 13184
rect 4212 13132 4218 13184
rect 4798 13132 4804 13184
rect 4856 13132 4862 13184
rect 6362 13132 6368 13184
rect 6420 13132 6426 13184
rect 6546 13132 6552 13184
rect 6604 13132 6610 13184
rect 6914 13132 6920 13184
rect 6972 13132 6978 13184
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 9125 13175 9183 13181
rect 9125 13172 9137 13175
rect 8812 13144 9137 13172
rect 8812 13132 8818 13144
rect 9125 13141 9137 13144
rect 9171 13141 9183 13175
rect 9232 13172 9260 13212
rect 9493 13209 9505 13243
rect 9539 13240 9551 13243
rect 9858 13240 9864 13252
rect 9539 13212 9864 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 11330 13200 11336 13252
rect 11388 13240 11394 13252
rect 11388 13212 14136 13240
rect 11388 13200 11394 13212
rect 9585 13175 9643 13181
rect 9585 13172 9597 13175
rect 9232 13144 9597 13172
rect 9125 13135 9183 13141
rect 9585 13141 9597 13144
rect 9631 13172 9643 13175
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9631 13144 10425 13172
rect 9631 13141 9643 13144
rect 9585 13135 9643 13141
rect 10413 13141 10425 13144
rect 10459 13172 10471 13175
rect 10502 13172 10508 13184
rect 10459 13144 10508 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11149 13175 11207 13181
rect 11149 13172 11161 13175
rect 11112 13144 11161 13172
rect 11112 13132 11118 13144
rect 11149 13141 11161 13144
rect 11195 13141 11207 13175
rect 11149 13135 11207 13141
rect 13078 13132 13084 13184
rect 13136 13132 13142 13184
rect 14108 13172 14136 13212
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14338 13243 14396 13249
rect 14338 13240 14350 13243
rect 14240 13212 14350 13240
rect 14240 13200 14246 13212
rect 14338 13209 14350 13212
rect 14384 13209 14396 13243
rect 14338 13203 14396 13209
rect 16592 13172 16620 13280
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 16942 13268 16948 13320
rect 17000 13268 17006 13320
rect 18046 13268 18052 13320
rect 18104 13308 18110 13320
rect 18892 13317 18920 13348
rect 22002 13336 22008 13388
rect 22060 13376 22066 13388
rect 24765 13379 24823 13385
rect 24765 13376 24777 13379
rect 22060 13348 24777 13376
rect 22060 13336 22066 13348
rect 24765 13345 24777 13348
rect 24811 13345 24823 13379
rect 24765 13339 24823 13345
rect 25038 13336 25044 13388
rect 25096 13336 25102 13388
rect 26234 13336 26240 13388
rect 26292 13336 26298 13388
rect 18509 13311 18567 13317
rect 18509 13308 18521 13311
rect 18104 13280 18521 13308
rect 18104 13268 18110 13280
rect 18509 13277 18521 13280
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 20625 13311 20683 13317
rect 20625 13277 20637 13311
rect 20671 13308 20683 13311
rect 20714 13308 20720 13320
rect 20671 13280 20720 13308
rect 20671 13277 20683 13280
rect 20625 13271 20683 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 23109 13311 23167 13317
rect 23109 13277 23121 13311
rect 23155 13308 23167 13311
rect 24118 13308 24124 13320
rect 23155 13280 24124 13308
rect 23155 13277 23167 13280
rect 23109 13271 23167 13277
rect 24118 13268 24124 13280
rect 24176 13268 24182 13320
rect 26252 13308 26280 13336
rect 26174 13280 26280 13308
rect 17282 13243 17340 13249
rect 17282 13240 17294 13243
rect 16684 13212 17294 13240
rect 16684 13181 16712 13212
rect 17282 13209 17294 13212
rect 17328 13209 17340 13243
rect 17282 13203 17340 13209
rect 18138 13200 18144 13252
rect 18196 13240 18202 13252
rect 18693 13243 18751 13249
rect 18693 13240 18705 13243
rect 18196 13212 18705 13240
rect 18196 13200 18202 13212
rect 18693 13209 18705 13212
rect 18739 13209 18751 13243
rect 18693 13203 18751 13209
rect 18785 13243 18843 13249
rect 18785 13209 18797 13243
rect 18831 13209 18843 13243
rect 18785 13203 18843 13209
rect 14108 13144 16620 13172
rect 16669 13175 16727 13181
rect 16669 13141 16681 13175
rect 16715 13141 16727 13175
rect 16669 13135 16727 13141
rect 16758 13132 16764 13184
rect 16816 13132 16822 13184
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 18506 13172 18512 13184
rect 18463 13144 18512 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 18506 13132 18512 13144
rect 18564 13172 18570 13184
rect 18800 13172 18828 13203
rect 19334 13200 19340 13252
rect 19392 13240 19398 13252
rect 20358 13243 20416 13249
rect 20358 13240 20370 13243
rect 19392 13212 20370 13240
rect 19392 13200 19398 13212
rect 20358 13209 20370 13212
rect 20404 13209 20416 13243
rect 20358 13203 20416 13209
rect 18564 13144 18828 13172
rect 18564 13132 18570 13144
rect 25774 13132 25780 13184
rect 25832 13172 25838 13184
rect 26513 13175 26571 13181
rect 26513 13172 26525 13175
rect 25832 13144 26525 13172
rect 25832 13132 25838 13144
rect 26513 13141 26525 13144
rect 26559 13141 26571 13175
rect 26513 13135 26571 13141
rect 1104 13082 26864 13104
rect 1104 13030 3658 13082
rect 3710 13030 3722 13082
rect 3774 13030 3786 13082
rect 3838 13030 3850 13082
rect 3902 13030 3914 13082
rect 3966 13030 3978 13082
rect 4030 13030 7658 13082
rect 7710 13030 7722 13082
rect 7774 13030 7786 13082
rect 7838 13030 7850 13082
rect 7902 13030 7914 13082
rect 7966 13030 7978 13082
rect 8030 13030 11658 13082
rect 11710 13030 11722 13082
rect 11774 13030 11786 13082
rect 11838 13030 11850 13082
rect 11902 13030 11914 13082
rect 11966 13030 11978 13082
rect 12030 13030 15658 13082
rect 15710 13030 15722 13082
rect 15774 13030 15786 13082
rect 15838 13030 15850 13082
rect 15902 13030 15914 13082
rect 15966 13030 15978 13082
rect 16030 13030 19658 13082
rect 19710 13030 19722 13082
rect 19774 13030 19786 13082
rect 19838 13030 19850 13082
rect 19902 13030 19914 13082
rect 19966 13030 19978 13082
rect 20030 13030 23658 13082
rect 23710 13030 23722 13082
rect 23774 13030 23786 13082
rect 23838 13030 23850 13082
rect 23902 13030 23914 13082
rect 23966 13030 23978 13082
rect 24030 13030 26864 13082
rect 1104 13008 26864 13030
rect 2038 12928 2044 12980
rect 2096 12928 2102 12980
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 3789 12971 3847 12977
rect 3789 12968 3801 12971
rect 3016 12940 3801 12968
rect 3016 12928 3022 12940
rect 3789 12937 3801 12940
rect 3835 12937 3847 12971
rect 3789 12931 3847 12937
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4798 12968 4804 12980
rect 4203 12940 4804 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 2584 12903 2642 12909
rect 2584 12869 2596 12903
rect 2630 12900 2642 12903
rect 2774 12900 2780 12912
rect 2630 12872 2780 12900
rect 2630 12869 2642 12872
rect 2584 12863 2642 12869
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 842 12792 848 12844
rect 900 12832 906 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 900 12804 1409 12832
rect 900 12792 906 12804
rect 1397 12801 1409 12804
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 2314 12724 2320 12776
rect 2372 12724 2378 12776
rect 3697 12699 3755 12705
rect 3697 12665 3709 12699
rect 3743 12696 3755 12699
rect 4172 12696 4200 12931
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 6178 12928 6184 12980
rect 6236 12928 6242 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 6288 12940 7757 12968
rect 4985 12903 5043 12909
rect 4985 12869 4997 12903
rect 5031 12900 5043 12903
rect 5534 12900 5540 12912
rect 5031 12872 5540 12900
rect 5031 12869 5043 12872
rect 4985 12863 5043 12869
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 5813 12903 5871 12909
rect 5813 12869 5825 12903
rect 5859 12900 5871 12903
rect 6288 12900 6316 12940
rect 7745 12937 7757 12940
rect 7791 12968 7803 12971
rect 9953 12971 10011 12977
rect 7791 12940 8340 12968
rect 7791 12937 7803 12940
rect 7745 12931 7803 12937
rect 5859 12872 6316 12900
rect 5859 12869 5871 12872
rect 5813 12863 5871 12869
rect 6362 12860 6368 12912
rect 6420 12900 6426 12912
rect 6610 12903 6668 12909
rect 6610 12900 6622 12903
rect 6420 12872 6622 12900
rect 6420 12860 6426 12872
rect 6610 12869 6622 12872
rect 6656 12869 6668 12903
rect 6610 12863 6668 12869
rect 6730 12860 6736 12912
rect 6788 12860 6794 12912
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 7374 12900 7380 12912
rect 6972 12872 7380 12900
rect 6972 12860 6978 12872
rect 7374 12860 7380 12872
rect 7432 12900 7438 12912
rect 8113 12903 8171 12909
rect 8113 12900 8125 12903
rect 7432 12872 8125 12900
rect 7432 12860 7438 12872
rect 8113 12869 8125 12872
rect 8159 12869 8171 12903
rect 8113 12863 8171 12869
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4724 12804 5089 12832
rect 4724 12776 4752 12804
rect 5077 12801 5089 12804
rect 5123 12832 5135 12835
rect 5442 12832 5448 12844
rect 5123 12804 5448 12832
rect 5123 12801 5135 12804
rect 5077 12795 5135 12801
rect 5442 12792 5448 12804
rect 5500 12832 5506 12844
rect 6748 12832 6776 12860
rect 5500 12804 5580 12832
rect 5500 12792 5506 12804
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 3743 12668 4200 12696
rect 3743 12665 3755 12668
rect 3697 12659 3755 12665
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 4264 12628 4292 12727
rect 4338 12724 4344 12776
rect 4396 12724 4402 12776
rect 4706 12724 4712 12776
rect 4764 12724 4770 12776
rect 5258 12724 5264 12776
rect 5316 12724 5322 12776
rect 4356 12696 4384 12724
rect 5442 12696 5448 12708
rect 4356 12668 5448 12696
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 5552 12696 5580 12804
rect 5644 12804 6776 12832
rect 5644 12776 5672 12804
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 8018 12832 8024 12844
rect 7708 12804 8024 12832
rect 7708 12792 7714 12804
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8205 12835 8263 12841
rect 8205 12801 8217 12835
rect 8251 12801 8263 12835
rect 8312 12832 8340 12940
rect 9953 12937 9965 12971
rect 9999 12968 10011 12971
rect 10686 12968 10692 12980
rect 9999 12940 10692 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11572 12940 11897 12968
rect 11572 12928 11578 12940
rect 11885 12937 11897 12940
rect 11931 12937 11943 12971
rect 11885 12931 11943 12937
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12253 12971 12311 12977
rect 12253 12968 12265 12971
rect 12216 12940 12265 12968
rect 12216 12928 12222 12940
rect 12253 12937 12265 12940
rect 12299 12937 12311 12971
rect 12253 12931 12311 12937
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14458 12968 14464 12980
rect 14415 12940 14464 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 15378 12968 15384 12980
rect 14783 12940 15384 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 16482 12928 16488 12980
rect 16540 12968 16546 12980
rect 16540 12940 17356 12968
rect 16540 12928 16546 12940
rect 9214 12860 9220 12912
rect 9272 12900 9278 12912
rect 12888 12903 12946 12909
rect 9272 12872 11652 12900
rect 9272 12860 9278 12872
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8312 12804 8401 12832
rect 8205 12795 8263 12801
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 5626 12724 5632 12776
rect 5684 12724 5690 12776
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5721 12727 5779 12733
rect 5736 12696 5764 12727
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 6365 12767 6423 12773
rect 6365 12764 6377 12767
rect 6052 12736 6377 12764
rect 6052 12724 6058 12736
rect 6365 12733 6377 12736
rect 6411 12733 6423 12767
rect 8220 12764 8248 12795
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 8737 12835 8795 12841
rect 8737 12832 8749 12835
rect 8628 12804 8749 12832
rect 8628 12792 8634 12804
rect 8737 12801 8749 12804
rect 8783 12801 8795 12835
rect 8737 12795 8795 12801
rect 9950 12792 9956 12844
rect 10008 12832 10014 12844
rect 10226 12832 10232 12844
rect 10008 12804 10232 12832
rect 10008 12792 10014 12804
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 11054 12792 11060 12844
rect 11112 12841 11118 12844
rect 11112 12832 11124 12841
rect 11112 12804 11157 12832
rect 11112 12795 11124 12804
rect 11112 12792 11118 12795
rect 8294 12764 8300 12776
rect 8220 12736 8300 12764
rect 6365 12727 6423 12733
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 8478 12724 8484 12776
rect 8536 12724 8542 12776
rect 11333 12767 11391 12773
rect 11333 12733 11345 12767
rect 11379 12733 11391 12767
rect 11333 12727 11391 12733
rect 5552 12668 5764 12696
rect 4120 12600 4292 12628
rect 4617 12631 4675 12637
rect 4120 12588 4126 12600
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 4798 12628 4804 12640
rect 4663 12600 4804 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 5736 12628 5764 12668
rect 7558 12656 7564 12708
rect 7616 12696 7622 12708
rect 7837 12699 7895 12705
rect 7837 12696 7849 12699
rect 7616 12668 7849 12696
rect 7616 12656 7622 12668
rect 7837 12665 7849 12668
rect 7883 12665 7895 12699
rect 11348 12696 11376 12727
rect 11514 12724 11520 12776
rect 11572 12764 11578 12776
rect 11624 12773 11652 12872
rect 12888 12869 12900 12903
rect 12934 12900 12946 12903
rect 13078 12900 13084 12912
rect 12934 12872 13084 12900
rect 12934 12869 12946 12872
rect 12888 12863 12946 12869
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 14826 12860 14832 12912
rect 14884 12860 14890 12912
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 16914 12903 16972 12909
rect 16914 12900 16926 12903
rect 16816 12872 16926 12900
rect 16816 12860 16822 12872
rect 16914 12869 16926 12872
rect 16960 12869 16972 12903
rect 17328 12900 17356 12940
rect 18046 12928 18052 12980
rect 18104 12928 18110 12980
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12937 18199 12971
rect 18141 12931 18199 12937
rect 18156 12900 18184 12931
rect 18506 12928 18512 12980
rect 18564 12928 18570 12980
rect 18601 12971 18659 12977
rect 18601 12937 18613 12971
rect 18647 12968 18659 12971
rect 18690 12968 18696 12980
rect 18647 12940 18696 12968
rect 18647 12937 18659 12940
rect 18601 12931 18659 12937
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 19242 12928 19248 12980
rect 19300 12968 19306 12980
rect 19337 12971 19395 12977
rect 19337 12968 19349 12971
rect 19300 12940 19349 12968
rect 19300 12928 19306 12940
rect 19337 12937 19349 12940
rect 19383 12937 19395 12971
rect 19337 12931 19395 12937
rect 19426 12928 19432 12980
rect 19484 12928 19490 12980
rect 19981 12971 20039 12977
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 20070 12968 20076 12980
rect 20027 12940 20076 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 24394 12928 24400 12980
rect 24452 12968 24458 12980
rect 24452 12940 26372 12968
rect 24452 12928 24458 12940
rect 17328 12872 18184 12900
rect 16914 12863 16972 12869
rect 19518 12860 19524 12912
rect 19576 12860 19582 12912
rect 26053 12903 26111 12909
rect 26053 12869 26065 12903
rect 26099 12900 26111 12903
rect 26142 12900 26148 12912
rect 26099 12872 26148 12900
rect 26099 12869 26111 12872
rect 26053 12863 26111 12869
rect 26142 12860 26148 12872
rect 26200 12860 26206 12912
rect 11716 12804 12434 12832
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11572 12736 11621 12764
rect 11572 12724 11578 12736
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 11716 12696 11744 12804
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 7837 12659 7895 12665
rect 9416 12668 10364 12696
rect 11348 12668 11744 12696
rect 9416 12628 9444 12668
rect 5736 12600 9444 12628
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 10226 12628 10232 12640
rect 9916 12600 10232 12628
rect 9916 12588 9922 12600
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 10336 12628 10364 12668
rect 11808 12628 11836 12727
rect 12406 12696 12434 12804
rect 14090 12792 14096 12844
rect 14148 12832 14154 12844
rect 19536 12832 19564 12860
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 14148 12804 18828 12832
rect 19536 12804 19809 12832
rect 14148 12792 14154 12804
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 12636 12696 12664 12727
rect 14918 12724 14924 12776
rect 14976 12724 14982 12776
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12733 16727 12767
rect 16669 12727 16727 12733
rect 12406 12668 12664 12696
rect 10336 12600 11836 12628
rect 12636 12628 12664 12668
rect 13556 12668 14872 12696
rect 13556 12628 13584 12668
rect 14844 12640 14872 12668
rect 12636 12600 13584 12628
rect 13998 12588 14004 12640
rect 14056 12588 14062 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 16684 12628 16712 12727
rect 18046 12724 18052 12776
rect 18104 12764 18110 12776
rect 18230 12764 18236 12776
rect 18104 12736 18236 12764
rect 18104 12724 18110 12736
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12733 18751 12767
rect 18800 12764 18828 12804
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 24946 12792 24952 12844
rect 25004 12792 25010 12844
rect 26344 12841 26372 12940
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 19426 12764 19432 12776
rect 18800 12736 19432 12764
rect 18693 12727 18751 12733
rect 17954 12656 17960 12708
rect 18012 12696 18018 12708
rect 18708 12696 18736 12727
rect 19426 12724 19432 12736
rect 19484 12764 19490 12776
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 19484 12736 19533 12764
rect 19484 12724 19490 12736
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 18012 12668 18736 12696
rect 18012 12656 18018 12668
rect 14884 12600 16712 12628
rect 14884 12588 14890 12600
rect 18782 12588 18788 12640
rect 18840 12628 18846 12640
rect 18969 12631 19027 12637
rect 18969 12628 18981 12631
rect 18840 12600 18981 12628
rect 18840 12588 18846 12600
rect 18969 12597 18981 12600
rect 19015 12597 19027 12631
rect 18969 12591 19027 12597
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 21821 12631 21879 12637
rect 21821 12628 21833 12631
rect 21232 12600 21833 12628
rect 21232 12588 21238 12600
rect 21821 12597 21833 12600
rect 21867 12597 21879 12631
rect 21821 12591 21879 12597
rect 24578 12588 24584 12640
rect 24636 12588 24642 12640
rect 1104 12538 26864 12560
rect 1104 12486 2918 12538
rect 2970 12486 2982 12538
rect 3034 12486 3046 12538
rect 3098 12486 3110 12538
rect 3162 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 6918 12538
rect 6970 12486 6982 12538
rect 7034 12486 7046 12538
rect 7098 12486 7110 12538
rect 7162 12486 7174 12538
rect 7226 12486 7238 12538
rect 7290 12486 10918 12538
rect 10970 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 11238 12538
rect 11290 12486 14918 12538
rect 14970 12486 14982 12538
rect 15034 12486 15046 12538
rect 15098 12486 15110 12538
rect 15162 12486 15174 12538
rect 15226 12486 15238 12538
rect 15290 12486 18918 12538
rect 18970 12486 18982 12538
rect 19034 12486 19046 12538
rect 19098 12486 19110 12538
rect 19162 12486 19174 12538
rect 19226 12486 19238 12538
rect 19290 12486 22918 12538
rect 22970 12486 22982 12538
rect 23034 12486 23046 12538
rect 23098 12486 23110 12538
rect 23162 12486 23174 12538
rect 23226 12486 23238 12538
rect 23290 12486 26864 12538
rect 1104 12464 26864 12486
rect 3237 12427 3295 12433
rect 3237 12393 3249 12427
rect 3283 12424 3295 12427
rect 4154 12424 4160 12436
rect 3283 12396 4160 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5534 12384 5540 12436
rect 5592 12384 5598 12436
rect 7374 12384 7380 12436
rect 7432 12384 7438 12436
rect 8570 12384 8576 12436
rect 8628 12384 8634 12436
rect 13081 12427 13139 12433
rect 13081 12393 13093 12427
rect 13127 12424 13139 12427
rect 13262 12424 13268 12436
rect 13127 12396 13268 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 18969 12427 19027 12433
rect 18969 12393 18981 12427
rect 19015 12424 19027 12427
rect 19334 12424 19340 12436
rect 19015 12396 19340 12424
rect 19015 12393 19027 12396
rect 18969 12387 19027 12393
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 22186 12384 22192 12436
rect 22244 12424 22250 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 22244 12396 22661 12424
rect 22244 12384 22250 12396
rect 22649 12393 22661 12396
rect 22695 12393 22707 12427
rect 22649 12387 22707 12393
rect 10042 12316 10048 12368
rect 10100 12356 10106 12368
rect 10100 12328 11100 12356
rect 10100 12316 10106 12328
rect 5994 12248 6000 12300
rect 6052 12248 6058 12300
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 8938 12288 8944 12300
rect 8536 12260 8944 12288
rect 8536 12248 8542 12260
rect 8938 12248 8944 12260
rect 8996 12288 9002 12300
rect 9033 12291 9091 12297
rect 9033 12288 9045 12291
rect 8996 12260 9045 12288
rect 8996 12248 9002 12260
rect 9033 12257 9045 12260
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 10502 12248 10508 12300
rect 10560 12288 10566 12300
rect 11072 12297 11100 12328
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 10560 12260 10977 12288
rect 10560 12248 10566 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11057 12291 11115 12297
rect 11057 12257 11069 12291
rect 11103 12257 11115 12291
rect 11057 12251 11115 12257
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 14734 12288 14740 12300
rect 13771 12260 14740 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20772 12260 20913 12288
rect 20772 12248 20778 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 21174 12248 21180 12300
rect 21232 12248 21238 12300
rect 24946 12248 24952 12300
rect 25004 12248 25010 12300
rect 1578 12180 1584 12232
rect 1636 12220 1642 12232
rect 1857 12223 1915 12229
rect 1857 12220 1869 12223
rect 1636 12192 1869 12220
rect 1636 12180 1642 12192
rect 1857 12189 1869 12192
rect 1903 12220 1915 12223
rect 1903 12192 2360 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 2332 12164 2360 12192
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 5534 12220 5540 12232
rect 4203 12192 5540 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 2130 12161 2136 12164
rect 2124 12152 2136 12161
rect 2091 12124 2136 12152
rect 2124 12115 2136 12124
rect 2130 12112 2136 12115
rect 2188 12112 2194 12164
rect 2314 12112 2320 12164
rect 2372 12152 2378 12164
rect 4172 12152 4200 12183
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 6012 12220 6040 12248
rect 5592 12192 6040 12220
rect 5592 12180 5598 12192
rect 8754 12180 8760 12232
rect 8812 12180 8818 12232
rect 18782 12180 18788 12232
rect 18840 12180 18846 12232
rect 20806 12180 20812 12232
rect 20864 12180 20870 12232
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 22925 12223 22983 12229
rect 22925 12220 22937 12223
rect 22796 12192 22937 12220
rect 22796 12180 22802 12192
rect 22925 12189 22937 12192
rect 22971 12189 22983 12223
rect 22925 12183 22983 12189
rect 23937 12223 23995 12229
rect 23937 12189 23949 12223
rect 23983 12220 23995 12223
rect 23983 12192 24440 12220
rect 23983 12189 23995 12192
rect 23937 12183 23995 12189
rect 2372 12124 4200 12152
rect 4424 12155 4482 12161
rect 2372 12112 2378 12124
rect 4424 12121 4436 12155
rect 4470 12152 4482 12155
rect 4614 12152 4620 12164
rect 4470 12124 4620 12152
rect 4470 12121 4482 12124
rect 4424 12115 4482 12121
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 6264 12155 6322 12161
rect 6264 12121 6276 12155
rect 6310 12152 6322 12155
rect 6362 12152 6368 12164
rect 6310 12124 6368 12152
rect 6310 12121 6322 12124
rect 6264 12115 6322 12121
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 9300 12155 9358 12161
rect 9300 12121 9312 12155
rect 9346 12152 9358 12155
rect 9398 12152 9404 12164
rect 9346 12124 9404 12152
rect 9346 12121 9358 12124
rect 9300 12115 9358 12121
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 10686 12152 10692 12164
rect 10428 12124 10692 12152
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4706 12084 4712 12096
rect 3927 12056 4712 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 10428 12093 10456 12124
rect 10686 12112 10692 12124
rect 10744 12152 10750 12164
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10744 12124 10885 12152
rect 10744 12112 10750 12124
rect 10873 12121 10885 12124
rect 10919 12121 10931 12155
rect 10873 12115 10931 12121
rect 13449 12155 13507 12161
rect 13449 12121 13461 12155
rect 13495 12152 13507 12155
rect 13998 12152 14004 12164
rect 13495 12124 14004 12152
rect 13495 12121 13507 12124
rect 13449 12115 13507 12121
rect 13998 12112 14004 12124
rect 14056 12112 14062 12164
rect 22833 12155 22891 12161
rect 22833 12152 22845 12155
rect 22402 12124 22845 12152
rect 22833 12121 22845 12124
rect 22879 12121 22891 12155
rect 22833 12115 22891 12121
rect 10413 12087 10471 12093
rect 10413 12053 10425 12087
rect 10459 12053 10471 12087
rect 10413 12047 10471 12053
rect 10502 12044 10508 12096
rect 10560 12044 10566 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13354 12084 13360 12096
rect 12952 12056 13360 12084
rect 12952 12044 12958 12056
rect 13354 12044 13360 12056
rect 13412 12084 13418 12096
rect 13541 12087 13599 12093
rect 13541 12084 13553 12087
rect 13412 12056 13553 12084
rect 13412 12044 13418 12056
rect 13541 12053 13553 12056
rect 13587 12053 13599 12087
rect 13541 12047 13599 12053
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20625 12087 20683 12093
rect 20625 12084 20637 12087
rect 20220 12056 20637 12084
rect 20220 12044 20226 12056
rect 20625 12053 20637 12056
rect 20671 12053 20683 12087
rect 20625 12047 20683 12053
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 24412 12093 24440 12192
rect 24762 12180 24768 12232
rect 24820 12180 24826 12232
rect 25774 12180 25780 12232
rect 25832 12180 25838 12232
rect 23753 12087 23811 12093
rect 23753 12084 23765 12087
rect 23624 12056 23765 12084
rect 23624 12044 23630 12056
rect 23753 12053 23765 12056
rect 23799 12053 23811 12087
rect 23753 12047 23811 12053
rect 24397 12087 24455 12093
rect 24397 12053 24409 12087
rect 24443 12053 24455 12087
rect 24397 12047 24455 12053
rect 24486 12044 24492 12096
rect 24544 12084 24550 12096
rect 24857 12087 24915 12093
rect 24857 12084 24869 12087
rect 24544 12056 24869 12084
rect 24544 12044 24550 12056
rect 24857 12053 24869 12056
rect 24903 12053 24915 12087
rect 24857 12047 24915 12053
rect 25685 12087 25743 12093
rect 25685 12053 25697 12087
rect 25731 12084 25743 12087
rect 25774 12084 25780 12096
rect 25731 12056 25780 12084
rect 25731 12053 25743 12056
rect 25685 12047 25743 12053
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 1104 11994 26864 12016
rect 1104 11942 3658 11994
rect 3710 11942 3722 11994
rect 3774 11942 3786 11994
rect 3838 11942 3850 11994
rect 3902 11942 3914 11994
rect 3966 11942 3978 11994
rect 4030 11942 7658 11994
rect 7710 11942 7722 11994
rect 7774 11942 7786 11994
rect 7838 11942 7850 11994
rect 7902 11942 7914 11994
rect 7966 11942 7978 11994
rect 8030 11942 11658 11994
rect 11710 11942 11722 11994
rect 11774 11942 11786 11994
rect 11838 11942 11850 11994
rect 11902 11942 11914 11994
rect 11966 11942 11978 11994
rect 12030 11942 15658 11994
rect 15710 11942 15722 11994
rect 15774 11942 15786 11994
rect 15838 11942 15850 11994
rect 15902 11942 15914 11994
rect 15966 11942 15978 11994
rect 16030 11942 19658 11994
rect 19710 11942 19722 11994
rect 19774 11942 19786 11994
rect 19838 11942 19850 11994
rect 19902 11942 19914 11994
rect 19966 11942 19978 11994
rect 20030 11942 23658 11994
rect 23710 11942 23722 11994
rect 23774 11942 23786 11994
rect 23838 11942 23850 11994
rect 23902 11942 23914 11994
rect 23966 11942 23978 11994
rect 24030 11942 26864 11994
rect 1104 11920 26864 11942
rect 2961 11883 3019 11889
rect 2961 11849 2973 11883
rect 3007 11880 3019 11883
rect 3007 11852 3464 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 1578 11704 1584 11756
rect 1636 11704 1642 11756
rect 1848 11747 1906 11753
rect 1848 11713 1860 11747
rect 1894 11744 1906 11747
rect 2130 11744 2136 11756
rect 1894 11716 2136 11744
rect 1894 11713 1906 11716
rect 1848 11707 1906 11713
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 3436 11753 3464 11852
rect 4614 11840 4620 11892
rect 4672 11840 4678 11892
rect 5902 11840 5908 11892
rect 5960 11840 5966 11892
rect 6362 11840 6368 11892
rect 6420 11840 6426 11892
rect 9398 11840 9404 11892
rect 9456 11840 9462 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9858 11880 9864 11892
rect 9732 11852 9864 11880
rect 9732 11840 9738 11852
rect 9858 11840 9864 11852
rect 9916 11880 9922 11892
rect 10965 11883 11023 11889
rect 9916 11852 10640 11880
rect 9916 11840 9922 11852
rect 10502 11812 10508 11824
rect 9600 11784 10508 11812
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11744 3479 11747
rect 4157 11747 4215 11753
rect 4157 11744 4169 11747
rect 3467 11716 4169 11744
rect 3467 11713 3479 11716
rect 3421 11707 3479 11713
rect 4157 11713 4169 11716
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4522 11744 4528 11756
rect 4387 11716 4528 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 4798 11704 4804 11756
rect 4856 11704 4862 11756
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 6086 11744 6092 11756
rect 5776 11716 6092 11744
rect 5776 11704 5782 11716
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6546 11704 6552 11756
rect 6604 11704 6610 11756
rect 9600 11753 9628 11784
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 10612 11821 10640 11852
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 12250 11880 12256 11892
rect 11011 11852 12256 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21637 11883 21695 11889
rect 21637 11880 21649 11883
rect 21048 11852 21649 11880
rect 21048 11840 21054 11852
rect 21637 11849 21649 11852
rect 21683 11849 21695 11883
rect 21637 11843 21695 11849
rect 22002 11840 22008 11892
rect 22060 11840 22066 11892
rect 22186 11840 22192 11892
rect 22244 11880 22250 11892
rect 22373 11883 22431 11889
rect 22373 11880 22385 11883
rect 22244 11852 22385 11880
rect 22244 11840 22250 11852
rect 22373 11849 22385 11852
rect 22419 11849 22431 11883
rect 22373 11843 22431 11849
rect 22738 11840 22744 11892
rect 22796 11880 22802 11892
rect 22796 11852 25452 11880
rect 22796 11840 22802 11852
rect 10597 11815 10655 11821
rect 10597 11781 10609 11815
rect 10643 11781 10655 11815
rect 10597 11775 10655 11781
rect 10686 11772 10692 11824
rect 10744 11772 10750 11824
rect 20162 11772 20168 11824
rect 20220 11772 20226 11824
rect 21726 11812 21732 11824
rect 21390 11784 21732 11812
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 23661 11815 23719 11821
rect 23661 11812 23673 11815
rect 23624 11784 23673 11812
rect 23624 11772 23630 11784
rect 23661 11781 23673 11784
rect 23707 11781 23719 11815
rect 25317 11815 25375 11821
rect 25317 11812 25329 11815
rect 24886 11784 25329 11812
rect 23661 11775 23719 11781
rect 25317 11781 25329 11784
rect 25363 11781 25375 11815
rect 25317 11775 25375 11781
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10376 11716 10425 11744
rect 10376 11704 10382 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 11330 11744 11336 11756
rect 10827 11716 11336 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 13998 11704 14004 11756
rect 14056 11704 14062 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 16666 11744 16672 11756
rect 14139 11716 16672 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 3384 11648 3525 11676
rect 3384 11636 3390 11648
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3694 11636 3700 11688
rect 3752 11636 3758 11688
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 14108 11676 14136 11707
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 25424 11753 25452 11852
rect 25409 11747 25467 11753
rect 25409 11713 25421 11747
rect 25455 11744 25467 11747
rect 25501 11747 25559 11753
rect 25501 11744 25513 11747
rect 25455 11716 25513 11744
rect 25455 11713 25467 11716
rect 25409 11707 25467 11713
rect 25501 11713 25513 11716
rect 25547 11713 25559 11747
rect 25501 11707 25559 11713
rect 9456 11648 14136 11676
rect 19889 11679 19947 11685
rect 9456 11636 9462 11648
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 21450 11676 21456 11688
rect 19935 11648 21456 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 21450 11636 21456 11648
rect 21508 11636 21514 11688
rect 22462 11636 22468 11688
rect 22520 11636 22526 11688
rect 22557 11679 22615 11685
rect 22557 11645 22569 11679
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 2590 11568 2596 11620
rect 2648 11608 2654 11620
rect 3053 11611 3111 11617
rect 3053 11608 3065 11611
rect 2648 11580 3065 11608
rect 2648 11568 2654 11580
rect 3053 11577 3065 11580
rect 3099 11577 3111 11611
rect 3053 11571 3111 11577
rect 21358 11568 21364 11620
rect 21416 11608 21422 11620
rect 22572 11608 22600 11639
rect 23382 11636 23388 11688
rect 23440 11636 23446 11688
rect 24946 11676 24952 11688
rect 23492 11648 24952 11676
rect 23492 11608 23520 11648
rect 24946 11636 24952 11648
rect 25004 11636 25010 11688
rect 21416 11580 23520 11608
rect 21416 11568 21422 11580
rect 24762 11568 24768 11620
rect 24820 11608 24826 11620
rect 25133 11611 25191 11617
rect 25133 11608 25145 11611
rect 24820 11580 25145 11608
rect 24820 11568 24826 11580
rect 25133 11577 25145 11580
rect 25179 11577 25191 11611
rect 25133 11571 25191 11577
rect 4525 11543 4583 11549
rect 4525 11509 4537 11543
rect 4571 11540 4583 11543
rect 6362 11540 6368 11552
rect 4571 11512 6368 11540
rect 4571 11509 4583 11512
rect 4525 11503 4583 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 14458 11540 14464 11552
rect 14323 11512 14464 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 25593 11543 25651 11549
rect 25593 11509 25605 11543
rect 25639 11540 25651 11543
rect 25682 11540 25688 11552
rect 25639 11512 25688 11540
rect 25639 11509 25651 11512
rect 25593 11503 25651 11509
rect 25682 11500 25688 11512
rect 25740 11500 25746 11552
rect 1104 11450 26864 11472
rect 1104 11398 2918 11450
rect 2970 11398 2982 11450
rect 3034 11398 3046 11450
rect 3098 11398 3110 11450
rect 3162 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 6918 11450
rect 6970 11398 6982 11450
rect 7034 11398 7046 11450
rect 7098 11398 7110 11450
rect 7162 11398 7174 11450
rect 7226 11398 7238 11450
rect 7290 11398 10918 11450
rect 10970 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 11238 11450
rect 11290 11398 14918 11450
rect 14970 11398 14982 11450
rect 15034 11398 15046 11450
rect 15098 11398 15110 11450
rect 15162 11398 15174 11450
rect 15226 11398 15238 11450
rect 15290 11398 18918 11450
rect 18970 11398 18982 11450
rect 19034 11398 19046 11450
rect 19098 11398 19110 11450
rect 19162 11398 19174 11450
rect 19226 11398 19238 11450
rect 19290 11398 22918 11450
rect 22970 11398 22982 11450
rect 23034 11398 23046 11450
rect 23098 11398 23110 11450
rect 23162 11398 23174 11450
rect 23226 11398 23238 11450
rect 23290 11398 26864 11450
rect 1104 11376 26864 11398
rect 2130 11296 2136 11348
rect 2188 11296 2194 11348
rect 12912 11308 17991 11336
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11237 12403 11271
rect 12345 11231 12403 11237
rect 8312 11172 9444 11200
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2590 11132 2596 11144
rect 2363 11104 2596 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2590 11092 2596 11104
rect 2648 11092 2654 11144
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8202 11132 8208 11144
rect 8067 11104 8208 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8312 11064 8340 11172
rect 9416 11144 9444 11172
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 7760 11036 8340 11064
rect 9048 11064 9076 11095
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 9306 11092 9312 11144
rect 9364 11092 9370 11144
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11132 12311 11135
rect 12360 11132 12388 11231
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 12912 11209 12940 11308
rect 15473 11271 15531 11277
rect 15473 11237 15485 11271
rect 15519 11237 15531 11271
rect 16298 11268 16304 11280
rect 15473 11231 15531 11237
rect 15948 11240 16304 11268
rect 12897 11203 12955 11209
rect 12897 11200 12909 11203
rect 12768 11172 12909 11200
rect 12768 11160 12774 11172
rect 12897 11169 12909 11172
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 12299 11104 12388 11132
rect 15381 11135 15439 11141
rect 12299 11101 12311 11104
rect 12253 11095 12311 11101
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15488 11132 15516 11231
rect 15948 11209 15976 11240
rect 16298 11228 16304 11240
rect 16356 11268 16362 11280
rect 16356 11240 17908 11268
rect 16356 11228 16362 11240
rect 15933 11203 15991 11209
rect 15933 11169 15945 11203
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 17770 11200 17776 11212
rect 16163 11172 17776 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16132 11132 16160 11163
rect 17770 11160 17776 11172
rect 17828 11160 17834 11212
rect 15427 11104 15516 11132
rect 15580 11104 16160 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 12158 11064 12164 11076
rect 9048 11036 12164 11064
rect 4154 10956 4160 11008
rect 4212 10996 4218 11008
rect 5166 10996 5172 11008
rect 4212 10968 5172 10996
rect 4212 10956 4218 10968
rect 5166 10956 5172 10968
rect 5224 10996 5230 11008
rect 7760 10996 7788 11036
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 14734 11064 14740 11076
rect 13228 11036 14740 11064
rect 13228 11024 13234 11036
rect 14734 11024 14740 11036
rect 14792 11064 14798 11076
rect 15580 11064 15608 11104
rect 14792 11036 15608 11064
rect 15841 11067 15899 11073
rect 14792 11024 14798 11036
rect 15841 11033 15853 11067
rect 15887 11064 15899 11067
rect 16298 11064 16304 11076
rect 15887 11036 16304 11064
rect 15887 11033 15899 11036
rect 15841 11027 15899 11033
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 5224 10968 7788 10996
rect 7837 10999 7895 11005
rect 5224 10956 5230 10968
rect 7837 10965 7849 10999
rect 7883 10996 7895 10999
rect 8110 10996 8116 11008
rect 7883 10968 8116 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 9582 10956 9588 11008
rect 9640 10956 9646 11008
rect 12066 10956 12072 11008
rect 12124 10956 12130 11008
rect 12710 10956 12716 11008
rect 12768 10956 12774 11008
rect 12805 10999 12863 11005
rect 12805 10965 12817 10999
rect 12851 10996 12863 10999
rect 12894 10996 12900 11008
rect 12851 10968 12900 10996
rect 12851 10965 12863 10968
rect 12805 10959 12863 10965
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 15194 10956 15200 11008
rect 15252 10956 15258 11008
rect 17880 10996 17908 11240
rect 17963 11200 17991 11308
rect 20806 11296 20812 11348
rect 20864 11296 20870 11348
rect 21726 11296 21732 11348
rect 21784 11296 21790 11348
rect 26050 11296 26056 11348
rect 26108 11336 26114 11348
rect 26145 11339 26203 11345
rect 26145 11336 26157 11339
rect 26108 11308 26157 11336
rect 26108 11296 26114 11308
rect 26145 11305 26157 11308
rect 26191 11305 26203 11339
rect 26145 11299 26203 11305
rect 18785 11271 18843 11277
rect 18785 11237 18797 11271
rect 18831 11268 18843 11271
rect 19518 11268 19524 11280
rect 18831 11240 19524 11268
rect 18831 11237 18843 11240
rect 18785 11231 18843 11237
rect 19518 11228 19524 11240
rect 19576 11228 19582 11280
rect 18141 11203 18199 11209
rect 18141 11200 18153 11203
rect 17963 11172 18153 11200
rect 18141 11169 18153 11172
rect 18187 11200 18199 11203
rect 18187 11172 19334 11200
rect 18187 11169 18199 11172
rect 18141 11163 18199 11169
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 19061 11135 19119 11141
rect 19061 11132 19073 11135
rect 18748 11104 19073 11132
rect 18748 11092 18754 11104
rect 19061 11101 19073 11104
rect 19107 11101 19119 11135
rect 19061 11095 19119 11101
rect 19306 11064 19334 11172
rect 21358 11160 21364 11212
rect 21416 11160 21422 11212
rect 21450 11160 21456 11212
rect 21508 11200 21514 11212
rect 23382 11200 23388 11212
rect 21508 11172 23388 11200
rect 21508 11160 21514 11172
rect 23382 11160 23388 11172
rect 23440 11200 23446 11212
rect 24397 11203 24455 11209
rect 24397 11200 24409 11203
rect 23440 11172 24409 11200
rect 23440 11160 23446 11172
rect 24397 11169 24409 11172
rect 24443 11169 24455 11203
rect 24397 11163 24455 11169
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 21048 11104 21189 11132
rect 21048 11092 21054 11104
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21821 11135 21879 11141
rect 21821 11101 21833 11135
rect 21867 11132 21879 11135
rect 22094 11132 22100 11144
rect 21867 11104 22100 11132
rect 21867 11101 21879 11104
rect 21821 11095 21879 11101
rect 22094 11092 22100 11104
rect 22152 11132 22158 11144
rect 22738 11132 22744 11144
rect 22152 11104 22744 11132
rect 22152 11092 22158 11104
rect 22738 11092 22744 11104
rect 22796 11132 22802 11144
rect 23569 11135 23627 11141
rect 23569 11132 23581 11135
rect 22796 11104 23581 11132
rect 22796 11092 22802 11104
rect 23569 11101 23581 11104
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 20162 11064 20168 11076
rect 19306 11036 20168 11064
rect 20162 11024 20168 11036
rect 20220 11064 20226 11076
rect 20438 11064 20444 11076
rect 20220 11036 20444 11064
rect 20220 11024 20226 11036
rect 20438 11024 20444 11036
rect 20496 11024 20502 11076
rect 21269 11067 21327 11073
rect 21269 11033 21281 11067
rect 21315 11064 21327 11067
rect 21542 11064 21548 11076
rect 21315 11036 21548 11064
rect 21315 11033 21327 11036
rect 21269 11027 21327 11033
rect 21542 11024 21548 11036
rect 21600 11024 21606 11076
rect 23845 11067 23903 11073
rect 23845 11033 23857 11067
rect 23891 11064 23903 11067
rect 24118 11064 24124 11076
rect 23891 11036 24124 11064
rect 23891 11033 23903 11036
rect 23845 11027 23903 11033
rect 24118 11024 24124 11036
rect 24176 11024 24182 11076
rect 24670 11024 24676 11076
rect 24728 11024 24734 11076
rect 25682 11024 25688 11076
rect 25740 11024 25746 11076
rect 18230 10996 18236 11008
rect 17880 10968 18236 10996
rect 18230 10956 18236 10968
rect 18288 10996 18294 11008
rect 18325 10999 18383 11005
rect 18325 10996 18337 10999
rect 18288 10968 18337 10996
rect 18288 10956 18294 10968
rect 18325 10965 18337 10968
rect 18371 10965 18383 10999
rect 18325 10959 18383 10965
rect 18414 10956 18420 11008
rect 18472 10956 18478 11008
rect 18874 10956 18880 11008
rect 18932 10956 18938 11008
rect 1104 10906 26864 10928
rect 1104 10854 3658 10906
rect 3710 10854 3722 10906
rect 3774 10854 3786 10906
rect 3838 10854 3850 10906
rect 3902 10854 3914 10906
rect 3966 10854 3978 10906
rect 4030 10854 7658 10906
rect 7710 10854 7722 10906
rect 7774 10854 7786 10906
rect 7838 10854 7850 10906
rect 7902 10854 7914 10906
rect 7966 10854 7978 10906
rect 8030 10854 11658 10906
rect 11710 10854 11722 10906
rect 11774 10854 11786 10906
rect 11838 10854 11850 10906
rect 11902 10854 11914 10906
rect 11966 10854 11978 10906
rect 12030 10854 15658 10906
rect 15710 10854 15722 10906
rect 15774 10854 15786 10906
rect 15838 10854 15850 10906
rect 15902 10854 15914 10906
rect 15966 10854 15978 10906
rect 16030 10854 19658 10906
rect 19710 10854 19722 10906
rect 19774 10854 19786 10906
rect 19838 10854 19850 10906
rect 19902 10854 19914 10906
rect 19966 10854 19978 10906
rect 20030 10854 23658 10906
rect 23710 10854 23722 10906
rect 23774 10854 23786 10906
rect 23838 10854 23850 10906
rect 23902 10854 23914 10906
rect 23966 10854 23978 10906
rect 24030 10854 26864 10906
rect 1104 10832 26864 10854
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10761 4399 10795
rect 4341 10755 4399 10761
rect 2774 10684 2780 10736
rect 2832 10724 2838 10736
rect 3418 10724 3424 10736
rect 2832 10696 3424 10724
rect 2832 10684 2838 10696
rect 3418 10684 3424 10696
rect 3476 10724 3482 10736
rect 4065 10727 4123 10733
rect 4065 10724 4077 10727
rect 3476 10696 4077 10724
rect 3476 10684 3482 10696
rect 4065 10693 4077 10696
rect 4111 10693 4123 10727
rect 4065 10687 4123 10693
rect 3786 10616 3792 10668
rect 3844 10616 3850 10668
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 1394 10548 1400 10600
rect 1452 10548 1458 10600
rect 3988 10588 4016 10619
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 4356 10656 4384 10755
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 7558 10792 7564 10804
rect 5040 10764 5212 10792
rect 5040 10752 5046 10764
rect 5184 10733 5212 10764
rect 6932 10764 7564 10792
rect 5169 10727 5227 10733
rect 5169 10693 5181 10727
rect 5215 10693 5227 10727
rect 5169 10687 5227 10693
rect 5074 10665 5080 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4356 10628 4905 10656
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5041 10659 5080 10665
rect 5041 10625 5053 10659
rect 5041 10619 5080 10625
rect 5074 10616 5080 10619
rect 5132 10616 5138 10668
rect 5258 10616 5264 10668
rect 5316 10616 5322 10668
rect 5350 10616 5356 10668
rect 5408 10665 5414 10668
rect 5408 10659 5457 10665
rect 5408 10625 5411 10659
rect 5445 10656 5457 10659
rect 6730 10656 6736 10668
rect 5445 10628 6736 10656
rect 5445 10625 5457 10628
rect 5408 10619 5457 10625
rect 5408 10616 5414 10619
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 6932 10665 6960 10764
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 7668 10764 9076 10792
rect 7009 10727 7067 10733
rect 7009 10693 7021 10727
rect 7055 10724 7067 10727
rect 7374 10724 7380 10736
rect 7055 10696 7380 10724
rect 7055 10693 7067 10696
rect 7009 10687 7067 10693
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 7668 10724 7696 10764
rect 8938 10724 8944 10736
rect 7484 10696 7696 10724
rect 7760 10696 8944 10724
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 4798 10588 4804 10600
rect 3988 10560 4804 10588
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 7116 10588 7144 10619
rect 7190 10616 7196 10668
rect 7248 10656 7254 10668
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 7248 10628 7297 10656
rect 7248 10616 7254 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7484 10588 7512 10696
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7760 10656 7788 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 9048 10724 9076 10764
rect 10042 10752 10048 10804
rect 10100 10752 10106 10804
rect 10134 10752 10140 10804
rect 10192 10752 10198 10804
rect 11422 10792 11428 10804
rect 10244 10764 11428 10792
rect 10244 10724 10272 10764
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 13170 10792 13176 10804
rect 11532 10764 13176 10792
rect 9048 10696 10272 10724
rect 7607 10628 7788 10656
rect 7828 10659 7886 10665
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7828 10625 7840 10659
rect 7874 10656 7886 10659
rect 8110 10656 8116 10668
rect 7874 10628 8116 10656
rect 7874 10625 7886 10628
rect 7828 10619 7886 10625
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 9456 10628 9505 10656
rect 9456 10616 9462 10628
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9582 10616 9588 10668
rect 9640 10616 9646 10668
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 7116 10560 7512 10588
rect 9784 10588 9812 10619
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 10313 10659 10371 10665
rect 10313 10656 10325 10659
rect 9916 10628 10325 10656
rect 9916 10616 9922 10628
rect 10313 10625 10325 10628
rect 10359 10625 10371 10659
rect 10313 10619 10371 10625
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10560 10628 10609 10656
rect 10560 10616 10566 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 10226 10588 10232 10600
rect 9784 10560 10232 10588
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 7190 10480 7196 10532
rect 7248 10520 7254 10532
rect 7466 10520 7472 10532
rect 7248 10492 7472 10520
rect 7248 10480 7254 10492
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 9490 10480 9496 10532
rect 9548 10520 9554 10532
rect 10704 10520 10732 10619
rect 9548 10492 10732 10520
rect 9548 10480 9554 10492
rect 1486 10412 1492 10464
rect 1544 10452 1550 10464
rect 2041 10455 2099 10461
rect 2041 10452 2053 10455
rect 1544 10424 2053 10452
rect 1544 10412 1550 10424
rect 2041 10421 2053 10424
rect 2087 10421 2099 10455
rect 2041 10415 2099 10421
rect 5537 10455 5595 10461
rect 5537 10421 5549 10455
rect 5583 10452 5595 10455
rect 5902 10452 5908 10464
rect 5583 10424 5908 10452
rect 5583 10421 5595 10424
rect 5537 10415 5595 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 6733 10455 6791 10461
rect 6733 10452 6745 10455
rect 6144 10424 6745 10452
rect 6144 10412 6150 10424
rect 6733 10421 6745 10424
rect 6779 10421 6791 10455
rect 6733 10415 6791 10421
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 8941 10455 8999 10461
rect 8941 10452 8953 10455
rect 8352 10424 8953 10452
rect 8352 10412 8358 10424
rect 8941 10421 8953 10424
rect 8987 10452 8999 10455
rect 9306 10452 9312 10464
rect 8987 10424 9312 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 11532 10452 11560 10764
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 13446 10792 13452 10804
rect 13311 10764 13452 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 13446 10752 13452 10764
rect 13504 10792 13510 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 13504 10764 13737 10792
rect 13504 10752 13510 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 13725 10755 13783 10761
rect 16298 10752 16304 10804
rect 16356 10752 16362 10804
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 17310 10792 17316 10804
rect 16816 10764 17316 10792
rect 16816 10752 16822 10764
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17589 10795 17647 10801
rect 17589 10761 17601 10795
rect 17635 10792 17647 10795
rect 17865 10795 17923 10801
rect 17865 10792 17877 10795
rect 17635 10764 17877 10792
rect 17635 10761 17647 10764
rect 17589 10755 17647 10761
rect 17865 10761 17877 10764
rect 17911 10792 17923 10795
rect 18414 10792 18420 10804
rect 17911 10764 18420 10792
rect 17911 10761 17923 10764
rect 17865 10755 17923 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10761 19395 10795
rect 19337 10755 19395 10761
rect 24305 10795 24363 10801
rect 24305 10761 24317 10795
rect 24351 10792 24363 10795
rect 24486 10792 24492 10804
rect 24351 10764 24492 10792
rect 24351 10761 24363 10764
rect 24305 10755 24363 10761
rect 15194 10733 15200 10736
rect 15188 10724 15200 10733
rect 11900 10696 14872 10724
rect 15155 10696 15200 10724
rect 11900 10665 11928 10696
rect 14844 10668 14872 10696
rect 15188 10687 15200 10696
rect 15194 10684 15200 10687
rect 15252 10684 15258 10736
rect 19000 10727 19058 10733
rect 19000 10693 19012 10727
rect 19046 10724 19058 10727
rect 19352 10724 19380 10755
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 24670 10752 24676 10804
rect 24728 10752 24734 10804
rect 25225 10795 25283 10801
rect 25225 10761 25237 10795
rect 25271 10792 25283 10795
rect 26050 10792 26056 10804
rect 25271 10764 26056 10792
rect 25271 10761 25283 10764
rect 25225 10755 25283 10761
rect 26050 10752 26056 10764
rect 26108 10752 26114 10804
rect 19046 10696 19380 10724
rect 20165 10727 20223 10733
rect 19046 10693 19058 10696
rect 19000 10687 19058 10693
rect 20165 10693 20177 10727
rect 20211 10724 20223 10727
rect 20254 10724 20260 10736
rect 20211 10696 20260 10724
rect 20211 10693 20223 10696
rect 20165 10687 20223 10693
rect 20254 10684 20260 10696
rect 20312 10684 20318 10736
rect 21910 10724 21916 10736
rect 21390 10696 21916 10724
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 25038 10724 25044 10736
rect 24412 10696 25044 10724
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 12141 10659 12199 10665
rect 12141 10656 12153 10659
rect 11885 10619 11943 10625
rect 11992 10628 12153 10656
rect 9640 10424 11560 10452
rect 11624 10452 11652 10619
rect 11992 10588 12020 10628
rect 12141 10625 12153 10628
rect 12187 10625 12199 10659
rect 12141 10619 12199 10625
rect 13170 10616 13176 10668
rect 13228 10656 13234 10668
rect 13722 10656 13728 10668
rect 13228 10628 13728 10656
rect 13228 10616 13234 10628
rect 13722 10616 13728 10628
rect 13780 10656 13786 10668
rect 13780 10628 13952 10656
rect 13780 10616 13786 10628
rect 11808 10560 12020 10588
rect 11808 10529 11836 10560
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 13924 10597 13952 10628
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 14056 10628 14197 10656
rect 14056 10616 14062 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14458 10616 14464 10668
rect 14516 10616 14522 10668
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14884 10628 14933 10656
rect 14884 10616 14890 10628
rect 14921 10625 14933 10628
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 17310 10616 17316 10668
rect 17368 10616 17374 10668
rect 17678 10616 17684 10668
rect 17736 10616 17742 10668
rect 19518 10616 19524 10668
rect 19576 10616 19582 10668
rect 24412 10665 24440 10696
rect 25038 10684 25044 10696
rect 25096 10684 25102 10736
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 24489 10659 24547 10665
rect 24489 10625 24501 10659
rect 24535 10656 24547 10659
rect 24535 10628 24900 10656
rect 24535 10625 24547 10628
rect 24489 10619 24547 10625
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 12952 10560 13829 10588
rect 12952 10548 12958 10560
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10588 14427 10591
rect 14734 10588 14740 10600
rect 14415 10560 14740 10588
rect 14415 10557 14427 10560
rect 14369 10551 14427 10557
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10588 19303 10591
rect 19889 10591 19947 10597
rect 19889 10588 19901 10591
rect 19291 10560 19901 10588
rect 19291 10557 19303 10560
rect 19245 10551 19303 10557
rect 19889 10557 19901 10560
rect 19935 10588 19947 10591
rect 21450 10588 21456 10600
rect 19935 10560 21456 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 24872 10529 24900 10628
rect 24946 10616 24952 10668
rect 25004 10656 25010 10668
rect 25004 10628 25452 10656
rect 25004 10616 25010 10628
rect 25424 10600 25452 10628
rect 25130 10548 25136 10600
rect 25188 10588 25194 10600
rect 25317 10591 25375 10597
rect 25317 10588 25329 10591
rect 25188 10560 25329 10588
rect 25188 10548 25194 10560
rect 25317 10557 25329 10560
rect 25363 10557 25375 10591
rect 25317 10551 25375 10557
rect 25406 10548 25412 10600
rect 25464 10548 25470 10600
rect 11793 10523 11851 10529
rect 11793 10489 11805 10523
rect 11839 10489 11851 10523
rect 13357 10523 13415 10529
rect 13357 10520 13369 10523
rect 11793 10483 11851 10489
rect 12912 10492 13369 10520
rect 12912 10452 12940 10492
rect 13357 10489 13369 10492
rect 13403 10489 13415 10523
rect 13357 10483 13415 10489
rect 24857 10523 24915 10529
rect 24857 10489 24869 10523
rect 24903 10489 24915 10523
rect 24857 10483 24915 10489
rect 11624 10424 12940 10452
rect 9640 10412 9646 10424
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14185 10455 14243 10461
rect 14185 10452 14197 10455
rect 13780 10424 14197 10452
rect 13780 10412 13786 10424
rect 14185 10421 14197 10424
rect 14231 10421 14243 10455
rect 14185 10415 14243 10421
rect 14642 10412 14648 10464
rect 14700 10412 14706 10464
rect 16942 10412 16948 10464
rect 17000 10412 17006 10464
rect 17218 10412 17224 10464
rect 17276 10412 17282 10464
rect 17402 10412 17408 10464
rect 17460 10412 17466 10464
rect 21637 10455 21695 10461
rect 21637 10421 21649 10455
rect 21683 10452 21695 10455
rect 21726 10452 21732 10464
rect 21683 10424 21732 10452
rect 21683 10421 21695 10424
rect 21637 10415 21695 10421
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 1104 10362 26864 10384
rect 1104 10310 2918 10362
rect 2970 10310 2982 10362
rect 3034 10310 3046 10362
rect 3098 10310 3110 10362
rect 3162 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 6918 10362
rect 6970 10310 6982 10362
rect 7034 10310 7046 10362
rect 7098 10310 7110 10362
rect 7162 10310 7174 10362
rect 7226 10310 7238 10362
rect 7290 10310 10918 10362
rect 10970 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 11238 10362
rect 11290 10310 14918 10362
rect 14970 10310 14982 10362
rect 15034 10310 15046 10362
rect 15098 10310 15110 10362
rect 15162 10310 15174 10362
rect 15226 10310 15238 10362
rect 15290 10310 18918 10362
rect 18970 10310 18982 10362
rect 19034 10310 19046 10362
rect 19098 10310 19110 10362
rect 19162 10310 19174 10362
rect 19226 10310 19238 10362
rect 19290 10310 22918 10362
rect 22970 10310 22982 10362
rect 23034 10310 23046 10362
rect 23098 10310 23110 10362
rect 23162 10310 23174 10362
rect 23226 10310 23238 10362
rect 23290 10310 26864 10362
rect 1104 10288 26864 10310
rect 3326 10248 3332 10260
rect 2746 10220 3332 10248
rect 2746 10180 2774 10220
rect 3326 10208 3332 10220
rect 3384 10248 3390 10260
rect 4522 10248 4528 10260
rect 3384 10220 4528 10248
rect 3384 10208 3390 10220
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 5408 10220 5672 10248
rect 5408 10208 5414 10220
rect 4154 10180 4160 10192
rect 2516 10152 2774 10180
rect 3528 10152 4160 10180
rect 2516 10121 2544 10152
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10081 2559 10115
rect 2501 10075 2559 10081
rect 2682 10072 2688 10124
rect 2740 10072 2746 10124
rect 3528 10121 3556 10152
rect 4154 10140 4160 10152
rect 4212 10180 4218 10192
rect 4430 10180 4436 10192
rect 4212 10152 4436 10180
rect 4212 10140 4218 10152
rect 4430 10140 4436 10152
rect 4488 10140 4494 10192
rect 5442 10180 5448 10192
rect 4540 10152 5448 10180
rect 3513 10115 3571 10121
rect 3513 10081 3525 10115
rect 3559 10081 3571 10115
rect 4540 10112 4568 10152
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 3513 10075 3571 10081
rect 3896 10084 4568 10112
rect 4709 10115 4767 10121
rect 1486 10004 1492 10056
rect 1544 10004 1550 10056
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 2774 10044 2780 10056
rect 2455 10016 2780 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3326 10044 3332 10056
rect 3283 10016 3332 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3326 10004 3332 10016
rect 3384 10044 3390 10056
rect 3786 10044 3792 10056
rect 3384 10016 3792 10044
rect 3384 10004 3390 10016
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 3896 9976 3924 10084
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 5166 10112 5172 10124
rect 4755 10084 5172 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 5166 10072 5172 10084
rect 5224 10112 5230 10124
rect 5644 10121 5672 10220
rect 6086 10208 6092 10260
rect 6144 10208 6150 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 7558 10248 7564 10260
rect 6319 10220 7564 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8202 10248 8208 10260
rect 7975 10220 8208 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 10318 10248 10324 10260
rect 8864 10220 10324 10248
rect 5994 10140 6000 10192
rect 6052 10180 6058 10192
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 6052 10152 6653 10180
rect 6052 10140 6058 10152
rect 6641 10149 6653 10152
rect 6687 10149 6699 10183
rect 6641 10143 6699 10149
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 6788 10152 7328 10180
rect 6788 10140 6794 10152
rect 5629 10115 5687 10121
rect 5224 10084 5488 10112
rect 5224 10072 5230 10084
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4019 10016 4108 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 1719 9948 3924 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 2041 9911 2099 9917
rect 2041 9908 2053 9911
rect 1912 9880 2053 9908
rect 1912 9868 1918 9880
rect 2041 9877 2053 9880
rect 2087 9877 2099 9911
rect 2041 9871 2099 9877
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 3344 9917 3372 9948
rect 2869 9911 2927 9917
rect 2869 9908 2881 9911
rect 2832 9880 2881 9908
rect 2832 9868 2838 9880
rect 2869 9877 2881 9880
rect 2915 9877 2927 9911
rect 2869 9871 2927 9877
rect 3329 9911 3387 9917
rect 3329 9877 3341 9911
rect 3375 9877 3387 9911
rect 3329 9871 3387 9877
rect 3789 9911 3847 9917
rect 3789 9877 3801 9911
rect 3835 9908 3847 9911
rect 3970 9908 3976 9920
rect 3835 9880 3976 9908
rect 3835 9877 3847 9880
rect 3789 9871 3847 9877
rect 3970 9868 3976 9880
rect 4028 9868 4034 9920
rect 4080 9917 4108 10016
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 5132 10016 5365 10044
rect 5132 10004 5138 10016
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 5258 9976 5264 9988
rect 4479 9948 5264 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 5460 9976 5488 10084
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 7098 10112 7104 10124
rect 5675 10084 7104 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 7190 10072 7196 10124
rect 7248 10072 7254 10124
rect 7300 10112 7328 10152
rect 7300 10084 8432 10112
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10044 6147 10047
rect 6362 10044 6368 10056
rect 6135 10016 6368 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 5368 9948 5488 9976
rect 5368 9920 5396 9948
rect 5810 9936 5816 9988
rect 5868 9936 5874 9988
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 6012 9976 6040 10007
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 7558 10044 7564 10056
rect 6595 10016 7564 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 8404 10044 8432 10084
rect 8478 10072 8484 10124
rect 8536 10072 8542 10124
rect 8570 10044 8576 10056
rect 8404 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8864 10044 8892 10220
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10468 10220 10701 10248
rect 10468 10208 10474 10220
rect 10689 10217 10701 10220
rect 10735 10217 10747 10251
rect 10689 10211 10747 10217
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12768 10220 13093 10248
rect 12768 10208 12774 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 13081 10211 13139 10217
rect 8938 10072 8944 10124
rect 8996 10112 9002 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8996 10084 9321 10112
rect 8996 10072 9002 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 8864 10016 9045 10044
rect 9033 10013 9045 10016
rect 9079 10013 9091 10047
rect 9324 10044 9352 10075
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 9324 10016 11713 10044
rect 9033 10007 9091 10013
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 13096 10044 13124 10211
rect 13722 10208 13728 10260
rect 13780 10208 13786 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16574 10248 16580 10260
rect 16448 10220 16580 10248
rect 16448 10208 16454 10220
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 17402 10248 17408 10260
rect 16899 10220 17408 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 17494 10208 17500 10260
rect 17552 10208 17558 10260
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 18874 10248 18880 10260
rect 17920 10220 18880 10248
rect 17920 10208 17926 10220
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 25130 10208 25136 10260
rect 25188 10208 25194 10260
rect 13372 10084 14780 10112
rect 13372 10053 13400 10084
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 13096 10016 13185 10044
rect 11701 10007 11759 10013
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14274 10044 14280 10056
rect 13872 10016 14280 10044
rect 13872 10004 13878 10016
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 7009 9979 7067 9985
rect 5960 9948 6040 9976
rect 6196 9948 6500 9976
rect 5960 9936 5966 9948
rect 4065 9911 4123 9917
rect 4065 9877 4077 9911
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 4522 9868 4528 9920
rect 4580 9868 4586 9920
rect 4982 9868 4988 9920
rect 5040 9868 5046 9920
rect 5350 9868 5356 9920
rect 5408 9868 5414 9920
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 6196 9908 6224 9948
rect 5500 9880 6224 9908
rect 5500 9868 5506 9880
rect 6362 9868 6368 9920
rect 6420 9868 6426 9920
rect 6472 9908 6500 9948
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 7374 9976 7380 9988
rect 7055 9948 7380 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 9554 9979 9612 9985
rect 9554 9976 9566 9979
rect 9232 9948 9566 9976
rect 7101 9911 7159 9917
rect 7101 9908 7113 9911
rect 6472 9880 7113 9908
rect 7101 9877 7113 9880
rect 7147 9908 7159 9911
rect 8110 9908 8116 9920
rect 7147 9880 8116 9908
rect 7147 9877 7159 9880
rect 7101 9871 7159 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 8662 9908 8668 9920
rect 8444 9880 8668 9908
rect 8444 9868 8450 9880
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 9232 9917 9260 9948
rect 9554 9945 9566 9948
rect 9600 9945 9612 9979
rect 9554 9939 9612 9945
rect 11968 9979 12026 9985
rect 11968 9945 11980 9979
rect 12014 9976 12026 9979
rect 12066 9976 12072 9988
rect 12014 9948 12072 9976
rect 12014 9945 12026 9948
rect 11968 9939 12026 9945
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 13630 9936 13636 9988
rect 13688 9976 13694 9988
rect 14384 9976 14412 10007
rect 14550 10004 14556 10056
rect 14608 10004 14614 10056
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 14752 10044 14780 10084
rect 14826 10072 14832 10124
rect 14884 10072 14890 10124
rect 17678 10112 17684 10124
rect 16132 10084 17684 10112
rect 16132 10044 16160 10084
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 19061 10115 19119 10121
rect 19061 10081 19073 10115
rect 19107 10112 19119 10115
rect 21450 10112 21456 10124
rect 19107 10084 21456 10112
rect 19107 10081 19119 10084
rect 19061 10075 19119 10081
rect 16301 10047 16359 10053
rect 16301 10044 16313 10047
rect 14752 10016 16160 10044
rect 16224 10016 16313 10044
rect 13688 9948 14412 9976
rect 15096 9979 15154 9985
rect 13688 9936 13694 9948
rect 15096 9945 15108 9979
rect 15142 9976 15154 9979
rect 15286 9976 15292 9988
rect 15142 9948 15292 9976
rect 15142 9945 15154 9948
rect 15096 9939 15154 9945
rect 15286 9936 15292 9948
rect 15344 9936 15350 9988
rect 16224 9920 16252 10016
rect 16301 10013 16313 10016
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16390 10004 16396 10056
rect 16448 10044 16454 10056
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 16448 10016 16589 10044
rect 16448 10004 16454 10016
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16666 10004 16672 10056
rect 16724 10004 16730 10056
rect 16942 10004 16948 10056
rect 17000 10004 17006 10056
rect 17034 10004 17040 10056
rect 17092 10004 17098 10056
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 17402 10044 17408 10056
rect 17359 10016 17408 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 16482 9936 16488 9988
rect 16540 9936 16546 9988
rect 17236 9976 17264 10007
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 19076 10044 19104 10075
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 21726 10072 21732 10124
rect 21784 10072 21790 10124
rect 18380 10016 19104 10044
rect 23477 10047 23535 10053
rect 18380 10004 18386 10016
rect 23477 10013 23489 10047
rect 23523 10044 23535 10047
rect 24118 10044 24124 10056
rect 23523 10016 24124 10044
rect 23523 10013 23535 10016
rect 23477 10007 23535 10013
rect 24118 10004 24124 10016
rect 24176 10044 24182 10056
rect 24762 10044 24768 10056
rect 24176 10016 24768 10044
rect 24176 10004 24182 10016
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 24854 10004 24860 10056
rect 24912 10004 24918 10056
rect 25038 10004 25044 10056
rect 25096 10004 25102 10056
rect 25222 10004 25228 10056
rect 25280 10044 25286 10056
rect 25317 10047 25375 10053
rect 25317 10044 25329 10047
rect 25280 10016 25329 10044
rect 25280 10004 25286 10016
rect 25317 10013 25329 10016
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 25501 10047 25559 10053
rect 25501 10013 25513 10047
rect 25547 10044 25559 10047
rect 25682 10044 25688 10056
rect 25547 10016 25688 10044
rect 25547 10013 25559 10016
rect 25501 10007 25559 10013
rect 25682 10004 25688 10016
rect 25740 10004 25746 10056
rect 26142 10004 26148 10056
rect 26200 10044 26206 10056
rect 26513 10047 26571 10053
rect 26513 10044 26525 10047
rect 26200 10016 26525 10044
rect 26200 10004 26206 10016
rect 26513 10013 26525 10016
rect 26559 10013 26571 10047
rect 26513 10007 26571 10013
rect 17236 9948 17724 9976
rect 9217 9911 9275 9917
rect 9217 9877 9229 9911
rect 9263 9877 9275 9911
rect 9217 9871 9275 9877
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 12492 9880 14105 9908
rect 12492 9868 12498 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 16206 9868 16212 9920
rect 16264 9868 16270 9920
rect 17696 9917 17724 9948
rect 18782 9936 18788 9988
rect 18840 9985 18846 9988
rect 18840 9976 18852 9985
rect 23385 9979 23443 9985
rect 23385 9976 23397 9979
rect 18840 9948 18885 9976
rect 22954 9948 23397 9976
rect 18840 9939 18852 9948
rect 23385 9945 23397 9948
rect 23431 9945 23443 9979
rect 23385 9939 23443 9945
rect 18840 9936 18846 9939
rect 17681 9911 17739 9917
rect 17681 9877 17693 9911
rect 17727 9908 17739 9911
rect 18414 9908 18420 9920
rect 17727 9880 18420 9908
rect 17727 9877 17739 9880
rect 17681 9871 17739 9877
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 23201 9911 23259 9917
rect 23201 9877 23213 9911
rect 23247 9908 23259 9911
rect 23290 9908 23296 9920
rect 23247 9880 23296 9908
rect 23247 9877 23259 9880
rect 23201 9871 23259 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 24946 9868 24952 9920
rect 25004 9868 25010 9920
rect 26326 9868 26332 9920
rect 26384 9868 26390 9920
rect 1104 9818 26864 9840
rect 1104 9766 3658 9818
rect 3710 9766 3722 9818
rect 3774 9766 3786 9818
rect 3838 9766 3850 9818
rect 3902 9766 3914 9818
rect 3966 9766 3978 9818
rect 4030 9766 7658 9818
rect 7710 9766 7722 9818
rect 7774 9766 7786 9818
rect 7838 9766 7850 9818
rect 7902 9766 7914 9818
rect 7966 9766 7978 9818
rect 8030 9766 11658 9818
rect 11710 9766 11722 9818
rect 11774 9766 11786 9818
rect 11838 9766 11850 9818
rect 11902 9766 11914 9818
rect 11966 9766 11978 9818
rect 12030 9766 15658 9818
rect 15710 9766 15722 9818
rect 15774 9766 15786 9818
rect 15838 9766 15850 9818
rect 15902 9766 15914 9818
rect 15966 9766 15978 9818
rect 16030 9766 19658 9818
rect 19710 9766 19722 9818
rect 19774 9766 19786 9818
rect 19838 9766 19850 9818
rect 19902 9766 19914 9818
rect 19966 9766 19978 9818
rect 20030 9766 23658 9818
rect 23710 9766 23722 9818
rect 23774 9766 23786 9818
rect 23838 9766 23850 9818
rect 23902 9766 23914 9818
rect 23966 9766 23978 9818
rect 24030 9766 26864 9818
rect 1104 9744 26864 9766
rect 3326 9664 3332 9716
rect 3384 9664 3390 9716
rect 4893 9707 4951 9713
rect 4893 9673 4905 9707
rect 4939 9704 4951 9707
rect 5258 9704 5264 9716
rect 4939 9676 5264 9704
rect 4939 9673 4951 9676
rect 4893 9667 4951 9673
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 6822 9704 6828 9716
rect 5408 9676 6828 9704
rect 5408 9664 5414 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7837 9707 7895 9713
rect 7837 9704 7849 9707
rect 7616 9676 7849 9704
rect 7616 9664 7622 9676
rect 7837 9673 7849 9676
rect 7883 9673 7895 9707
rect 7837 9667 7895 9673
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 10134 9704 10140 9716
rect 8168 9676 10140 9704
rect 8168 9664 8174 9676
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 10468 9676 10885 9704
rect 10468 9664 10474 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 10873 9667 10931 9673
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 14645 9707 14703 9713
rect 14645 9704 14657 9707
rect 14608 9676 14657 9704
rect 14608 9664 14614 9676
rect 14645 9673 14657 9676
rect 14691 9673 14703 9707
rect 14645 9667 14703 9673
rect 15286 9664 15292 9716
rect 15344 9664 15350 9716
rect 15933 9707 15991 9713
rect 15933 9673 15945 9707
rect 15979 9704 15991 9707
rect 16206 9704 16212 9716
rect 15979 9676 16212 9704
rect 15979 9673 15991 9676
rect 15933 9667 15991 9673
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 17034 9664 17040 9716
rect 17092 9704 17098 9716
rect 17681 9707 17739 9713
rect 17681 9704 17693 9707
rect 17092 9676 17693 9704
rect 17092 9664 17098 9676
rect 17681 9673 17693 9676
rect 17727 9673 17739 9707
rect 17681 9667 17739 9673
rect 18414 9664 18420 9716
rect 18472 9664 18478 9716
rect 24780 9676 25084 9704
rect 5534 9636 5540 9648
rect 1964 9608 5540 9636
rect 1854 9528 1860 9580
rect 1912 9528 1918 9580
rect 1964 9577 1992 9608
rect 3528 9580 3556 9608
rect 5534 9596 5540 9608
rect 5592 9636 5598 9648
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 5592 9608 5733 9636
rect 5592 9596 5598 9608
rect 5721 9605 5733 9608
rect 5767 9636 5779 9639
rect 5767 9608 6408 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2216 9571 2274 9577
rect 2216 9537 2228 9571
rect 2262 9568 2274 9571
rect 2682 9568 2688 9580
rect 2262 9540 2688 9568
rect 2262 9537 2274 9540
rect 2216 9531 2274 9537
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 1964 9500 1992 9531
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 3780 9571 3838 9577
rect 3568 9540 3593 9568
rect 3568 9528 3574 9540
rect 3780 9537 3792 9571
rect 3826 9568 3838 9571
rect 4062 9568 4068 9580
rect 3826 9540 4068 9568
rect 3826 9537 3838 9540
rect 3780 9531 3838 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5166 9568 5172 9580
rect 5031 9540 5172 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6380 9577 6408 9608
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 7524 9608 8217 9636
rect 7524 9596 7530 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 10229 9639 10287 9645
rect 10229 9636 10241 9639
rect 8205 9599 8263 9605
rect 8956 9608 10241 9636
rect 8956 9580 8984 9608
rect 10229 9605 10241 9608
rect 10275 9605 10287 9639
rect 10229 9599 10287 9605
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 12216 9608 17264 9636
rect 12216 9596 12222 9608
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 6621 9571 6679 9577
rect 6621 9568 6633 9571
rect 6365 9531 6423 9537
rect 6472 9540 6633 9568
rect 6472 9500 6500 9540
rect 6621 9537 6633 9540
rect 6667 9537 6679 9571
rect 6621 9531 6679 9537
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 7432 9540 7788 9568
rect 7432 9528 7438 9540
rect 1544 9472 1992 9500
rect 6196 9472 6500 9500
rect 1544 9460 1550 9472
rect 6196 9441 6224 9472
rect 6181 9435 6239 9441
rect 6181 9401 6193 9435
rect 6227 9401 6239 9435
rect 6181 9395 6239 9401
rect 1670 9324 1676 9376
rect 1728 9324 1734 9376
rect 7760 9373 7788 9540
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 8352 9540 8616 9568
rect 8352 9528 8358 9540
rect 8481 9503 8539 9509
rect 8481 9469 8493 9503
rect 8527 9469 8539 9503
rect 8588 9500 8616 9540
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 10594 9568 10600 9580
rect 9539 9540 10600 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 14108 9577 14136 9608
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 14182 9528 14188 9580
rect 14240 9528 14246 9580
rect 14366 9528 14372 9580
rect 14424 9528 14430 9580
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9537 14519 9571
rect 14461 9531 14519 9537
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9568 15531 9571
rect 16025 9571 16083 9577
rect 15519 9540 15608 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 9214 9500 9220 9512
rect 8588 9472 9220 9500
rect 8481 9463 8539 9469
rect 7745 9367 7803 9373
rect 7745 9333 7757 9367
rect 7791 9333 7803 9367
rect 8496 9364 8524 9463
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 10134 9460 10140 9512
rect 10192 9500 10198 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10192 9472 10977 9500
rect 10192 9460 10198 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11057 9503 11115 9509
rect 11057 9469 11069 9503
rect 11103 9500 11115 9503
rect 13446 9500 13452 9512
rect 11103 9472 13452 9500
rect 11103 9469 11115 9472
rect 11057 9463 11115 9469
rect 10318 9392 10324 9444
rect 10376 9432 10382 9444
rect 10505 9435 10563 9441
rect 10505 9432 10517 9435
rect 10376 9404 10517 9432
rect 10376 9392 10382 9404
rect 10505 9401 10517 9404
rect 10551 9401 10563 9435
rect 10505 9395 10563 9401
rect 10686 9392 10692 9444
rect 10744 9432 10750 9444
rect 11072 9432 11100 9463
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 10744 9404 11100 9432
rect 10744 9392 10750 9404
rect 11330 9392 11336 9444
rect 11388 9432 11394 9444
rect 11388 9404 11560 9432
rect 11388 9392 11394 9404
rect 11422 9364 11428 9376
rect 8496 9336 11428 9364
rect 7745 9327 7803 9333
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 11532 9364 11560 9404
rect 14476 9364 14504 9531
rect 15580 9441 15608 9540
rect 16025 9537 16037 9571
rect 16071 9568 16083 9571
rect 16390 9568 16396 9580
rect 16071 9540 16396 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 17236 9577 17264 9608
rect 18230 9596 18236 9648
rect 18288 9636 18294 9648
rect 18325 9639 18383 9645
rect 18325 9636 18337 9639
rect 18288 9608 18337 9636
rect 18288 9596 18294 9608
rect 18325 9605 18337 9608
rect 18371 9605 18383 9639
rect 18325 9599 18383 9605
rect 21910 9596 21916 9648
rect 21968 9596 21974 9648
rect 24780 9636 24808 9676
rect 22020 9608 24808 9636
rect 24923 9639 24981 9645
rect 17221 9571 17279 9577
rect 17221 9537 17233 9571
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 17586 9568 17592 9580
rect 17543 9540 17592 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 17773 9571 17831 9577
rect 17773 9537 17785 9571
rect 17819 9568 17831 9571
rect 17862 9568 17868 9580
rect 17819 9540 17868 9568
rect 17819 9537 17831 9540
rect 17773 9531 17831 9537
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 18414 9568 18420 9580
rect 18104 9540 18420 9568
rect 18104 9528 18110 9540
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 22020 9577 22048 9608
rect 24923 9605 24935 9639
rect 24969 9636 24981 9639
rect 25056 9636 25084 9676
rect 26326 9636 26332 9648
rect 24969 9605 24992 9636
rect 25056 9608 26332 9636
rect 24923 9599 24992 9605
rect 21637 9571 21695 9577
rect 21637 9537 21649 9571
rect 21683 9568 21695 9571
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21683 9540 22017 9568
rect 21683 9537 21695 9540
rect 21637 9531 21695 9537
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22830 9528 22836 9580
rect 22888 9568 22894 9580
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 22888 9540 23121 9568
rect 22888 9528 22894 9540
rect 23109 9537 23121 9540
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 24578 9528 24584 9580
rect 24636 9568 24642 9580
rect 24673 9571 24731 9577
rect 24673 9568 24685 9571
rect 24636 9540 24685 9568
rect 24636 9528 24642 9540
rect 24673 9537 24685 9540
rect 24719 9568 24731 9571
rect 24765 9571 24823 9577
rect 24765 9568 24777 9571
rect 24719 9540 24777 9568
rect 24719 9537 24731 9540
rect 24673 9531 24731 9537
rect 24765 9537 24777 9540
rect 24811 9537 24823 9571
rect 24765 9531 24823 9537
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9500 16267 9503
rect 16850 9500 16856 9512
rect 16255 9472 16856 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9500 18291 9503
rect 19334 9500 19340 9512
rect 18279 9472 19340 9500
rect 18279 9469 18291 9472
rect 18233 9463 18291 9469
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 21453 9503 21511 9509
rect 21453 9469 21465 9503
rect 21499 9469 21511 9503
rect 21453 9463 21511 9469
rect 15565 9435 15623 9441
rect 15565 9401 15577 9435
rect 15611 9401 15623 9435
rect 15565 9395 15623 9401
rect 18690 9392 18696 9444
rect 18748 9432 18754 9444
rect 18785 9435 18843 9441
rect 18785 9432 18797 9435
rect 18748 9404 18797 9432
rect 18748 9392 18754 9404
rect 18785 9401 18797 9404
rect 18831 9401 18843 9435
rect 18785 9395 18843 9401
rect 17494 9364 17500 9376
rect 11532 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17957 9367 18015 9373
rect 17957 9333 17969 9367
rect 18003 9364 18015 9367
rect 18046 9364 18052 9376
rect 18003 9336 18052 9364
rect 18003 9333 18015 9336
rect 17957 9327 18015 9333
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 21468 9364 21496 9463
rect 22462 9460 22468 9512
rect 22520 9500 22526 9512
rect 22741 9503 22799 9509
rect 22741 9500 22753 9503
rect 22520 9472 22753 9500
rect 22520 9460 22526 9472
rect 22741 9469 22753 9472
rect 22787 9469 22799 9503
rect 22741 9463 22799 9469
rect 23201 9503 23259 9509
rect 23201 9469 23213 9503
rect 23247 9500 23259 9503
rect 24210 9500 24216 9512
rect 23247 9472 24216 9500
rect 23247 9469 23259 9472
rect 23201 9463 23259 9469
rect 22756 9432 22784 9463
rect 24210 9460 24216 9472
rect 24268 9460 24274 9512
rect 24964 9432 24992 9599
rect 26326 9596 26332 9608
rect 26384 9596 26390 9648
rect 25041 9571 25099 9577
rect 25041 9537 25053 9571
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 25133 9571 25191 9577
rect 25133 9537 25145 9571
rect 25179 9537 25191 9571
rect 25133 9531 25191 9537
rect 22756 9404 24992 9432
rect 25056 9432 25084 9531
rect 25148 9500 25176 9531
rect 25222 9528 25228 9580
rect 25280 9568 25286 9580
rect 25501 9571 25559 9577
rect 25501 9568 25513 9571
rect 25280 9540 25513 9568
rect 25280 9528 25286 9540
rect 25501 9537 25513 9540
rect 25547 9537 25559 9571
rect 25501 9531 25559 9537
rect 25593 9571 25651 9577
rect 25593 9537 25605 9571
rect 25639 9568 25651 9571
rect 25682 9568 25688 9580
rect 25639 9540 25688 9568
rect 25639 9537 25651 9540
rect 25593 9531 25651 9537
rect 25608 9500 25636 9531
rect 25682 9528 25688 9540
rect 25740 9528 25746 9580
rect 25774 9528 25780 9580
rect 25832 9528 25838 9580
rect 25148 9472 25636 9500
rect 25792 9432 25820 9528
rect 25056 9404 25820 9432
rect 22094 9364 22100 9376
rect 21468 9336 22100 9364
rect 22094 9324 22100 9336
rect 22152 9364 22158 9376
rect 22646 9364 22652 9376
rect 22152 9336 22652 9364
rect 22152 9324 22158 9336
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23934 9324 23940 9376
rect 23992 9364 23998 9376
rect 24581 9367 24639 9373
rect 24581 9364 24593 9367
rect 23992 9336 24593 9364
rect 23992 9324 23998 9336
rect 24581 9333 24593 9336
rect 24627 9333 24639 9367
rect 24581 9327 24639 9333
rect 25409 9367 25467 9373
rect 25409 9333 25421 9367
rect 25455 9364 25467 9367
rect 25590 9364 25596 9376
rect 25455 9336 25596 9364
rect 25455 9333 25467 9336
rect 25409 9327 25467 9333
rect 25590 9324 25596 9336
rect 25648 9324 25654 9376
rect 25774 9324 25780 9376
rect 25832 9324 25838 9376
rect 1104 9274 26864 9296
rect 1104 9222 2918 9274
rect 2970 9222 2982 9274
rect 3034 9222 3046 9274
rect 3098 9222 3110 9274
rect 3162 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 6918 9274
rect 6970 9222 6982 9274
rect 7034 9222 7046 9274
rect 7098 9222 7110 9274
rect 7162 9222 7174 9274
rect 7226 9222 7238 9274
rect 7290 9222 10918 9274
rect 10970 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 11238 9274
rect 11290 9222 14918 9274
rect 14970 9222 14982 9274
rect 15034 9222 15046 9274
rect 15098 9222 15110 9274
rect 15162 9222 15174 9274
rect 15226 9222 15238 9274
rect 15290 9222 18918 9274
rect 18970 9222 18982 9274
rect 19034 9222 19046 9274
rect 19098 9222 19110 9274
rect 19162 9222 19174 9274
rect 19226 9222 19238 9274
rect 19290 9222 22918 9274
rect 22970 9222 22982 9274
rect 23034 9222 23046 9274
rect 23098 9222 23110 9274
rect 23162 9222 23174 9274
rect 23226 9222 23238 9274
rect 23290 9222 26864 9274
rect 1104 9200 26864 9222
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2740 9132 2973 9160
rect 2740 9120 2746 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 5132 9132 5181 9160
rect 5132 9120 5138 9132
rect 5169 9129 5181 9132
rect 5215 9129 5227 9163
rect 5169 9123 5227 9129
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7466 9160 7472 9172
rect 7331 9132 7472 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 13541 9163 13599 9169
rect 12492 9132 13492 9160
rect 12492 9120 12498 9132
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9092 2927 9095
rect 3418 9092 3424 9104
rect 2915 9064 3424 9092
rect 2915 9061 2927 9064
rect 2869 9055 2927 9061
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 13464 9092 13492 9132
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 14182 9160 14188 9172
rect 13587 9132 14188 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 16945 9163 17003 9169
rect 16945 9129 16957 9163
rect 16991 9160 17003 9163
rect 17402 9160 17408 9172
rect 16991 9132 17408 9160
rect 16991 9129 17003 9132
rect 16945 9123 17003 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 18104 9132 18460 9160
rect 18104 9120 18110 9132
rect 16482 9092 16488 9104
rect 9732 9064 13400 9092
rect 13464 9064 16488 9092
rect 9732 9052 9738 9064
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 3789 9027 3847 9033
rect 3789 9024 3801 9027
rect 3568 8996 3801 9024
rect 3568 8984 3574 8996
rect 3789 8993 3801 8996
rect 3835 8993 3847 9027
rect 3789 8987 3847 8993
rect 9214 8984 9220 9036
rect 9272 9024 9278 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 9272 8996 11161 9024
rect 9272 8984 9278 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 9024 11391 9027
rect 11379 8996 12572 9024
rect 11379 8993 11391 8996
rect 11333 8987 11391 8993
rect 1486 8916 1492 8968
rect 1544 8916 1550 8968
rect 1756 8959 1814 8965
rect 1756 8925 1768 8959
rect 1802 8925 1814 8959
rect 1756 8919 1814 8925
rect 1670 8848 1676 8900
rect 1728 8888 1734 8900
rect 1780 8888 1808 8919
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 3145 8959 3203 8965
rect 3145 8956 3157 8959
rect 2832 8928 3157 8956
rect 2832 8916 2838 8928
rect 3145 8925 3157 8928
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 4982 8956 4988 8968
rect 3467 8928 4988 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5592 8928 5733 8956
rect 5592 8916 5598 8928
rect 5721 8925 5733 8928
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 5902 8916 5908 8968
rect 5960 8916 5966 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9548 8928 9781 8956
rect 9548 8916 9554 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 4034 8891 4092 8897
rect 4034 8888 4046 8891
rect 1728 8860 1808 8888
rect 3620 8860 4046 8888
rect 1728 8848 1734 8860
rect 3620 8829 3648 8860
rect 4034 8857 4046 8860
rect 4080 8857 4092 8891
rect 4034 8851 4092 8857
rect 6172 8891 6230 8897
rect 6172 8857 6184 8891
rect 6218 8888 6230 8891
rect 6362 8888 6368 8900
rect 6218 8860 6368 8888
rect 6218 8857 6230 8860
rect 6172 8851 6230 8857
rect 6362 8848 6368 8860
rect 6420 8848 6426 8900
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8789 3663 8823
rect 3605 8783 3663 8789
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 8812 8792 10701 8820
rect 8812 8780 8818 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 10689 8783 10747 8789
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10836 8792 11069 8820
rect 10836 8780 10842 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 12434 8820 12440 8832
rect 11480 8792 12440 8820
rect 11480 8780 11486 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 12544 8820 12572 8996
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 13372 8965 13400 9064
rect 16482 9052 16488 9064
rect 16540 9052 16546 9104
rect 18322 8984 18328 9036
rect 18380 8984 18386 9036
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12676 8928 13001 8956
rect 12676 8916 12682 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12860 8860 13185 8888
rect 12860 8848 12866 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 13262 8848 13268 8900
rect 13320 8848 13326 8900
rect 13372 8888 13400 8919
rect 14826 8916 14832 8968
rect 14884 8916 14890 8968
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 17310 8956 17316 8968
rect 15436 8928 17316 8956
rect 15436 8916 15442 8928
rect 17310 8916 17316 8928
rect 17368 8916 17374 8968
rect 18058 8959 18116 8965
rect 18058 8925 18070 8959
rect 18104 8956 18116 8959
rect 18432 8956 18460 9132
rect 23566 9120 23572 9172
rect 23624 9160 23630 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 23624 9132 24409 9160
rect 23624 9120 23630 9132
rect 24397 9129 24409 9132
rect 24443 9129 24455 9163
rect 24397 9123 24455 9129
rect 24946 9120 24952 9172
rect 25004 9160 25010 9172
rect 25317 9163 25375 9169
rect 25317 9160 25329 9163
rect 25004 9132 25329 9160
rect 25004 9120 25010 9132
rect 25317 9129 25329 9132
rect 25363 9129 25375 9163
rect 25317 9123 25375 9129
rect 23477 9095 23535 9101
rect 23477 9061 23489 9095
rect 23523 9061 23535 9095
rect 23477 9055 23535 9061
rect 24213 9095 24271 9101
rect 24213 9061 24225 9095
rect 24259 9092 24271 9095
rect 24259 9064 25084 9092
rect 24259 9061 24271 9064
rect 24213 9055 24271 9061
rect 21450 8984 21456 9036
rect 21508 8984 21514 9036
rect 23201 9027 23259 9033
rect 23201 8993 23213 9027
rect 23247 9024 23259 9027
rect 23382 9024 23388 9036
rect 23247 8996 23388 9024
rect 23247 8993 23259 8996
rect 23201 8987 23259 8993
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 18104 8928 18460 8956
rect 18104 8925 18116 8928
rect 18058 8919 18116 8925
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 22554 8956 22560 8968
rect 21692 8928 22560 8956
rect 21692 8916 21698 8928
rect 22554 8916 22560 8928
rect 22612 8956 22618 8968
rect 23109 8959 23167 8965
rect 23109 8956 23121 8959
rect 22612 8928 23121 8956
rect 22612 8916 22618 8928
rect 23109 8925 23121 8928
rect 23155 8925 23167 8959
rect 23492 8956 23520 9055
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 23860 8996 24593 9024
rect 23569 8959 23627 8965
rect 23569 8956 23581 8959
rect 23492 8928 23581 8956
rect 23109 8919 23167 8925
rect 23569 8925 23581 8928
rect 23615 8925 23627 8959
rect 23569 8919 23627 8925
rect 23658 8916 23664 8968
rect 23716 8956 23722 8968
rect 23860 8956 23888 8996
rect 24581 8993 24593 8996
rect 24627 8993 24639 9027
rect 24581 8987 24639 8993
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 24949 9027 25007 9033
rect 24949 9024 24961 9027
rect 24912 8996 24961 9024
rect 24912 8984 24918 8996
rect 24949 8993 24961 8996
rect 24995 8993 25007 9027
rect 25056 9024 25084 9064
rect 25130 9052 25136 9104
rect 25188 9052 25194 9104
rect 25774 9024 25780 9036
rect 25056 8996 25268 9024
rect 24949 8987 25007 8993
rect 23716 8928 23888 8956
rect 23716 8916 23722 8928
rect 23934 8916 23940 8968
rect 23992 8916 23998 8968
rect 24118 8965 24124 8968
rect 24075 8959 24124 8965
rect 24075 8925 24087 8959
rect 24121 8925 24124 8959
rect 24075 8919 24124 8925
rect 24118 8916 24124 8919
rect 24176 8916 24182 8968
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 16574 8888 16580 8900
rect 13372 8860 16580 8888
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 20714 8848 20720 8900
rect 20772 8848 20778 8900
rect 21266 8848 21272 8900
rect 21324 8888 21330 8900
rect 21913 8891 21971 8897
rect 21913 8888 21925 8891
rect 21324 8860 21925 8888
rect 21324 8848 21330 8860
rect 21913 8857 21925 8860
rect 21959 8857 21971 8891
rect 21913 8851 21971 8857
rect 22281 8891 22339 8897
rect 22281 8857 22293 8891
rect 22327 8888 22339 8891
rect 23474 8888 23480 8900
rect 22327 8860 23480 8888
rect 22327 8857 22339 8860
rect 22281 8851 22339 8857
rect 23474 8848 23480 8860
rect 23532 8848 23538 8900
rect 23845 8891 23903 8897
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24688 8888 24716 8919
rect 24762 8916 24768 8968
rect 24820 8956 24826 8968
rect 24820 8928 25176 8956
rect 24820 8916 24826 8928
rect 23891 8860 24716 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 13814 8820 13820 8832
rect 12544 8792 13820 8820
rect 13814 8780 13820 8792
rect 13872 8820 13878 8832
rect 14550 8820 14556 8832
rect 13872 8792 14556 8820
rect 13872 8780 13878 8792
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 16482 8780 16488 8832
rect 16540 8820 16546 8832
rect 17954 8820 17960 8832
rect 16540 8792 17960 8820
rect 16540 8780 16546 8792
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 23566 8780 23572 8832
rect 23624 8820 23630 8832
rect 23860 8820 23888 8851
rect 24946 8848 24952 8900
rect 25004 8888 25010 8900
rect 25041 8891 25099 8897
rect 25041 8888 25053 8891
rect 25004 8860 25053 8888
rect 25004 8848 25010 8860
rect 25041 8857 25053 8860
rect 25087 8857 25099 8891
rect 25041 8851 25099 8857
rect 23624 8792 23888 8820
rect 25148 8820 25176 8928
rect 25240 8888 25268 8996
rect 25332 8996 25780 9024
rect 25332 8965 25360 8996
rect 25774 8984 25780 8996
rect 25832 8984 25838 9036
rect 25317 8959 25375 8965
rect 25317 8925 25329 8959
rect 25363 8925 25375 8959
rect 25317 8919 25375 8925
rect 25409 8959 25467 8965
rect 25409 8925 25421 8959
rect 25455 8925 25467 8959
rect 25409 8919 25467 8925
rect 25424 8888 25452 8919
rect 25590 8916 25596 8968
rect 25648 8916 25654 8968
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 25884 8888 25912 8919
rect 25240 8860 25452 8888
rect 25516 8860 25912 8888
rect 25516 8820 25544 8860
rect 25148 8792 25544 8820
rect 23624 8780 23630 8792
rect 25774 8780 25780 8832
rect 25832 8780 25838 8832
rect 1104 8730 26864 8752
rect 1104 8678 3658 8730
rect 3710 8678 3722 8730
rect 3774 8678 3786 8730
rect 3838 8678 3850 8730
rect 3902 8678 3914 8730
rect 3966 8678 3978 8730
rect 4030 8678 7658 8730
rect 7710 8678 7722 8730
rect 7774 8678 7786 8730
rect 7838 8678 7850 8730
rect 7902 8678 7914 8730
rect 7966 8678 7978 8730
rect 8030 8678 11658 8730
rect 11710 8678 11722 8730
rect 11774 8678 11786 8730
rect 11838 8678 11850 8730
rect 11902 8678 11914 8730
rect 11966 8678 11978 8730
rect 12030 8678 15658 8730
rect 15710 8678 15722 8730
rect 15774 8678 15786 8730
rect 15838 8678 15850 8730
rect 15902 8678 15914 8730
rect 15966 8678 15978 8730
rect 16030 8678 19658 8730
rect 19710 8678 19722 8730
rect 19774 8678 19786 8730
rect 19838 8678 19850 8730
rect 19902 8678 19914 8730
rect 19966 8678 19978 8730
rect 20030 8678 23658 8730
rect 23710 8678 23722 8730
rect 23774 8678 23786 8730
rect 23838 8678 23850 8730
rect 23902 8678 23914 8730
rect 23966 8678 23978 8730
rect 24030 8678 26864 8730
rect 1104 8656 26864 8678
rect 8941 8619 8999 8625
rect 8941 8585 8953 8619
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 5166 8508 5172 8560
rect 5224 8508 5230 8560
rect 8956 8548 8984 8579
rect 10502 8576 10508 8628
rect 10560 8576 10566 8628
rect 13814 8616 13820 8628
rect 12912 8588 13820 8616
rect 9278 8551 9336 8557
rect 9278 8548 9290 8551
rect 8956 8520 9290 8548
rect 9278 8517 9290 8520
rect 9324 8517 9336 8551
rect 12802 8548 12808 8560
rect 9278 8511 9336 8517
rect 10704 8520 12808 8548
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7374 8480 7380 8492
rect 7331 8452 7380 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 4908 8412 4936 8443
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 10704 8489 10732 8520
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8996 8452 9045 8480
rect 8996 8440 9002 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8480 11115 8483
rect 12158 8480 12164 8492
rect 11103 8452 12164 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 5902 8412 5908 8424
rect 4908 8384 5908 8412
rect 5902 8372 5908 8384
rect 5960 8412 5966 8424
rect 5997 8415 6055 8421
rect 5997 8412 6009 8415
rect 5960 8384 6009 8412
rect 5960 8372 5966 8384
rect 5997 8381 6009 8384
rect 6043 8412 6055 8415
rect 6454 8412 6460 8424
rect 6043 8384 6460 8412
rect 6043 8381 6055 8384
rect 5997 8375 6055 8381
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 10413 8347 10471 8353
rect 10413 8313 10425 8347
rect 10459 8344 10471 8347
rect 10796 8344 10824 8440
rect 10980 8412 11008 8443
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 11422 8412 11428 8424
rect 10980 8384 11428 8412
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 12710 8372 12716 8424
rect 12768 8372 12774 8424
rect 12912 8421 12940 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 14461 8619 14519 8625
rect 14461 8616 14473 8619
rect 14424 8588 14473 8616
rect 14424 8576 14430 8588
rect 14461 8585 14473 8588
rect 14507 8585 14519 8619
rect 14461 8579 14519 8585
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 14608 8588 15424 8616
rect 14608 8576 14614 8588
rect 14826 8548 14832 8560
rect 13096 8520 14832 8548
rect 13096 8489 13124 8520
rect 14826 8508 14832 8520
rect 14884 8548 14890 8560
rect 15289 8551 15347 8557
rect 15289 8548 15301 8551
rect 14884 8520 15301 8548
rect 14884 8508 14890 8520
rect 15289 8517 15301 8520
rect 15335 8517 15347 8551
rect 15396 8548 15424 8588
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17460 8588 17509 8616
rect 17460 8576 17466 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 17862 8576 17868 8628
rect 17920 8576 17926 8628
rect 20530 8616 20536 8628
rect 18800 8588 20536 8616
rect 18693 8551 18751 8557
rect 18693 8548 18705 8551
rect 15396 8520 18705 8548
rect 15289 8511 15347 8517
rect 18693 8517 18705 8520
rect 18739 8517 18751 8551
rect 18693 8511 18751 8517
rect 13354 8489 13360 8492
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13348 8443 13360 8489
rect 13354 8440 13360 8443
rect 13412 8440 13418 8492
rect 14550 8440 14556 8492
rect 14608 8440 14614 8492
rect 15746 8440 15752 8492
rect 15804 8440 15810 8492
rect 16390 8440 16396 8492
rect 16448 8480 16454 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 16448 8452 17417 8480
rect 16448 8440 16454 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8381 12955 8415
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 12897 8375 12955 8381
rect 14108 8384 17325 8412
rect 14108 8344 14136 8384
rect 17313 8381 17325 8384
rect 17359 8412 17371 8415
rect 18800 8412 18828 8588
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 21542 8616 21548 8628
rect 20640 8588 21548 8616
rect 20640 8557 20668 8588
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 23661 8619 23719 8625
rect 23661 8585 23673 8619
rect 23707 8616 23719 8619
rect 24118 8616 24124 8628
rect 23707 8588 24124 8616
rect 23707 8585 23719 8588
rect 23661 8579 23719 8585
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 20441 8551 20499 8557
rect 20441 8517 20453 8551
rect 20487 8517 20499 8551
rect 20441 8511 20499 8517
rect 20625 8551 20683 8557
rect 20625 8517 20637 8551
rect 20671 8517 20683 8551
rect 21910 8548 21916 8560
rect 20625 8511 20683 8517
rect 20732 8520 21916 8548
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 19705 8483 19763 8489
rect 19291 8452 19656 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 17359 8384 18828 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 19426 8372 19432 8424
rect 19484 8372 19490 8424
rect 19628 8412 19656 8452
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 20456 8480 20484 8511
rect 20732 8480 20760 8520
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 22465 8551 22523 8557
rect 22465 8548 22477 8551
rect 22296 8520 22477 8548
rect 19751 8452 20392 8480
rect 20456 8452 20760 8480
rect 21269 8483 21327 8489
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 19794 8412 19800 8424
rect 19628 8384 19800 8412
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 19889 8415 19947 8421
rect 19889 8381 19901 8415
rect 19935 8412 19947 8415
rect 19978 8412 19984 8424
rect 19935 8384 19984 8412
rect 19935 8381 19947 8384
rect 19889 8375 19947 8381
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 20162 8412 20168 8424
rect 20119 8384 20168 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20364 8412 20392 8452
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21450 8480 21456 8492
rect 21315 8452 21456 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 22296 8489 22324 8520
rect 22465 8517 22477 8520
rect 22511 8548 22523 8551
rect 25130 8548 25136 8560
rect 22511 8520 25136 8548
rect 22511 8517 22523 8520
rect 22465 8511 22523 8517
rect 25130 8508 25136 8520
rect 25188 8508 25194 8560
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 22830 8440 22836 8492
rect 22888 8480 22894 8492
rect 23293 8483 23351 8489
rect 23293 8480 23305 8483
rect 22888 8452 23305 8480
rect 22888 8440 22894 8452
rect 23293 8449 23305 8452
rect 23339 8449 23351 8483
rect 23293 8443 23351 8449
rect 21082 8412 21088 8424
rect 20364 8384 21088 8412
rect 21082 8372 21088 8384
rect 21140 8372 21146 8424
rect 21818 8372 21824 8424
rect 21876 8412 21882 8424
rect 22005 8415 22063 8421
rect 22005 8412 22017 8415
rect 21876 8384 22017 8412
rect 21876 8372 21882 8384
rect 22005 8381 22017 8384
rect 22051 8381 22063 8415
rect 22005 8375 22063 8381
rect 23385 8415 23443 8421
rect 23385 8381 23397 8415
rect 23431 8412 23443 8415
rect 24118 8412 24124 8424
rect 23431 8384 24124 8412
rect 23431 8381 23443 8384
rect 23385 8375 23443 8381
rect 24118 8372 24124 8384
rect 24176 8372 24182 8424
rect 10459 8316 10824 8344
rect 14016 8316 14136 8344
rect 10459 8313 10471 8316
rect 10413 8307 10471 8313
rect 7101 8279 7159 8285
rect 7101 8245 7113 8279
rect 7147 8276 7159 8279
rect 7466 8276 7472 8288
rect 7147 8248 7472 8276
rect 7147 8245 7159 8248
rect 7101 8239 7159 8245
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 12253 8279 12311 8285
rect 12253 8276 12265 8279
rect 11756 8248 12265 8276
rect 11756 8236 11762 8248
rect 12253 8245 12265 8248
rect 12299 8245 12311 8279
rect 12253 8239 12311 8245
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 14016 8276 14044 8316
rect 14550 8304 14556 8356
rect 14608 8344 14614 8356
rect 14608 8316 15240 8344
rect 14608 8304 14614 8316
rect 13504 8248 14044 8276
rect 15212 8276 15240 8316
rect 15562 8304 15568 8356
rect 15620 8304 15626 8356
rect 20257 8347 20315 8353
rect 20257 8313 20269 8347
rect 20303 8344 20315 8347
rect 20530 8344 20536 8356
rect 20303 8316 20536 8344
rect 20303 8313 20315 8316
rect 20257 8307 20315 8313
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 20714 8304 20720 8356
rect 20772 8344 20778 8356
rect 20772 8316 22094 8344
rect 20772 8304 20778 8316
rect 15470 8276 15476 8288
rect 15212 8248 15476 8276
rect 13504 8236 13510 8248
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 18598 8276 18604 8288
rect 15712 8248 18604 8276
rect 15712 8236 15718 8248
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 20441 8279 20499 8285
rect 20441 8245 20453 8279
rect 20487 8276 20499 8279
rect 21358 8276 21364 8288
rect 20487 8248 21364 8276
rect 20487 8245 20499 8248
rect 20441 8239 20499 8245
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 22066 8276 22094 8316
rect 22186 8276 22192 8288
rect 22066 8248 22192 8276
rect 22186 8236 22192 8248
rect 22244 8236 22250 8288
rect 22738 8236 22744 8288
rect 22796 8236 22802 8288
rect 1104 8186 26864 8208
rect 1104 8134 2918 8186
rect 2970 8134 2982 8186
rect 3034 8134 3046 8186
rect 3098 8134 3110 8186
rect 3162 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 6918 8186
rect 6970 8134 6982 8186
rect 7034 8134 7046 8186
rect 7098 8134 7110 8186
rect 7162 8134 7174 8186
rect 7226 8134 7238 8186
rect 7290 8134 10918 8186
rect 10970 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 11238 8186
rect 11290 8134 14918 8186
rect 14970 8134 14982 8186
rect 15034 8134 15046 8186
rect 15098 8134 15110 8186
rect 15162 8134 15174 8186
rect 15226 8134 15238 8186
rect 15290 8134 18918 8186
rect 18970 8134 18982 8186
rect 19034 8134 19046 8186
rect 19098 8134 19110 8186
rect 19162 8134 19174 8186
rect 19226 8134 19238 8186
rect 19290 8134 22918 8186
rect 22970 8134 22982 8186
rect 23034 8134 23046 8186
rect 23098 8134 23110 8186
rect 23162 8134 23174 8186
rect 23226 8134 23238 8186
rect 23290 8134 26864 8186
rect 1104 8112 26864 8134
rect 11422 8032 11428 8084
rect 11480 8032 11486 8084
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 12066 8072 12072 8084
rect 11747 8044 12072 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13412 8044 13553 8072
rect 13412 8032 13418 8044
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 15654 8072 15660 8084
rect 14700 8044 15660 8072
rect 14700 8032 14706 8044
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 15804 8044 15945 8072
rect 15804 8032 15810 8044
rect 15933 8041 15945 8044
rect 15979 8041 15991 8075
rect 15933 8035 15991 8041
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17184 8044 17325 8072
rect 17184 8032 17190 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 18230 8072 18236 8084
rect 17644 8044 18236 8072
rect 17644 8032 17650 8044
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 20809 8075 20867 8081
rect 20809 8072 20821 8075
rect 20772 8044 20821 8072
rect 20772 8032 20778 8044
rect 20809 8041 20821 8044
rect 20855 8041 20867 8075
rect 20809 8035 20867 8041
rect 23566 8032 23572 8084
rect 23624 8072 23630 8084
rect 23753 8075 23811 8081
rect 23753 8072 23765 8075
rect 23624 8044 23765 8072
rect 23624 8032 23630 8044
rect 23753 8041 23765 8044
rect 23799 8041 23811 8075
rect 23753 8035 23811 8041
rect 13449 8007 13507 8013
rect 13449 7973 13461 8007
rect 13495 8004 13507 8007
rect 13630 8004 13636 8016
rect 13495 7976 13636 8004
rect 13495 7973 13507 7976
rect 13449 7967 13507 7973
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 19337 8007 19395 8013
rect 13780 7976 14596 8004
rect 13780 7964 13786 7976
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 8996 7908 9413 7936
rect 8996 7896 9002 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 11422 7936 11428 7948
rect 9401 7899 9459 7905
rect 11072 7908 11428 7936
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6512 7840 6745 7868
rect 6512 7828 6518 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 7000 7871 7058 7877
rect 7000 7837 7012 7871
rect 7046 7868 7058 7871
rect 7466 7868 7472 7880
rect 7046 7840 7472 7868
rect 7046 7837 7058 7840
rect 7000 7831 7058 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 11072 7877 11100 7908
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 11606 7896 11612 7948
rect 11664 7936 11670 7948
rect 14568 7945 14596 7976
rect 16408 7976 17448 8004
rect 16408 7948 16436 7976
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11664 7908 12081 7936
rect 11664 7896 11670 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 14553 7939 14611 7945
rect 14553 7905 14565 7939
rect 14599 7905 14611 7939
rect 14553 7899 14611 7905
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 9232 7840 10885 7868
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 5534 7800 5540 7812
rect 4120 7772 5540 7800
rect 4120 7760 4126 7772
rect 5534 7760 5540 7772
rect 5592 7800 5598 7812
rect 8202 7800 8208 7812
rect 5592 7772 8208 7800
rect 5592 7760 5598 7772
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 9232 7732 9260 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7868 11299 7871
rect 11330 7868 11336 7880
rect 11287 7840 11336 7868
rect 11287 7837 11299 7840
rect 11241 7831 11299 7837
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 11698 7868 11704 7880
rect 11563 7840 11704 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 13262 7868 13268 7880
rect 11839 7840 13268 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 13771 7840 14136 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 9646 7803 9704 7809
rect 9646 7800 9658 7803
rect 9324 7772 9658 7800
rect 9324 7741 9352 7772
rect 9646 7769 9658 7772
rect 9692 7769 9704 7803
rect 9646 7763 9704 7769
rect 11149 7803 11207 7809
rect 11149 7769 11161 7803
rect 11195 7769 11207 7803
rect 12314 7803 12372 7809
rect 12314 7800 12326 7803
rect 11149 7763 11207 7769
rect 11992 7772 12326 7800
rect 8168 7704 9260 7732
rect 9309 7735 9367 7741
rect 8168 7692 8174 7704
rect 9309 7701 9321 7735
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11164 7732 11192 7763
rect 11992 7741 12020 7772
rect 12314 7769 12326 7772
rect 12360 7769 12372 7803
rect 12314 7763 12372 7769
rect 14108 7741 14136 7840
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14424 7840 14473 7868
rect 14424 7828 14430 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14660 7868 14688 7899
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 16390 7936 16396 7948
rect 16172 7908 16396 7936
rect 16172 7896 16178 7908
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16482 7896 16488 7948
rect 16540 7896 16546 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 16632 7908 17172 7936
rect 16632 7896 16638 7908
rect 14461 7831 14519 7837
rect 14568 7840 14688 7868
rect 14568 7812 14596 7840
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15528 7840 15853 7868
rect 15528 7828 15534 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 17144 7877 17172 7908
rect 17420 7877 17448 7976
rect 19337 7973 19349 8007
rect 19383 8004 19395 8007
rect 19702 8004 19708 8016
rect 19383 7976 19708 8004
rect 19383 7973 19395 7976
rect 19337 7967 19395 7973
rect 19702 7964 19708 7976
rect 19760 7964 19766 8016
rect 20162 7964 20168 8016
rect 20220 8004 20226 8016
rect 20220 7976 20668 8004
rect 20220 7964 20226 7976
rect 20640 7945 20668 7976
rect 20625 7939 20683 7945
rect 20625 7905 20637 7939
rect 20671 7905 20683 7939
rect 20625 7899 20683 7905
rect 21453 7939 21511 7945
rect 21453 7905 21465 7939
rect 21499 7936 21511 7939
rect 21818 7936 21824 7948
rect 21499 7908 21824 7936
rect 21499 7905 21511 7908
rect 21453 7899 21511 7905
rect 21818 7896 21824 7908
rect 21876 7896 21882 7948
rect 21910 7896 21916 7948
rect 21968 7896 21974 7948
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7936 22155 7939
rect 23290 7936 23296 7948
rect 22143 7908 23296 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 25958 7896 25964 7948
rect 26016 7936 26022 7948
rect 26513 7939 26571 7945
rect 26513 7936 26525 7939
rect 26016 7908 26525 7936
rect 26016 7896 26022 7908
rect 26513 7905 26525 7908
rect 26559 7905 26571 7939
rect 26513 7899 26571 7905
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16868 7840 17049 7868
rect 14182 7760 14188 7812
rect 14240 7800 14246 7812
rect 14550 7800 14556 7812
rect 14240 7772 14556 7800
rect 14240 7760 14246 7772
rect 14550 7760 14556 7772
rect 14608 7760 14614 7812
rect 14826 7760 14832 7812
rect 14884 7800 14890 7812
rect 15013 7803 15071 7809
rect 15013 7800 15025 7803
rect 14884 7772 15025 7800
rect 14884 7760 14890 7772
rect 15013 7769 15025 7772
rect 15059 7769 15071 7803
rect 15013 7763 15071 7769
rect 16301 7803 16359 7809
rect 16301 7769 16313 7803
rect 16347 7800 16359 7803
rect 16574 7800 16580 7812
rect 16347 7772 16580 7800
rect 16347 7769 16359 7772
rect 16301 7763 16359 7769
rect 16574 7760 16580 7772
rect 16632 7800 16638 7812
rect 16868 7800 16896 7840
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19484 7840 19717 7868
rect 19484 7828 19490 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19794 7828 19800 7880
rect 19852 7828 19858 7880
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 20128 7840 20177 7868
rect 20128 7828 20134 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 20530 7868 20536 7880
rect 20303 7840 20536 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 21174 7828 21180 7880
rect 21232 7868 21238 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 21232 7840 21281 7868
rect 21232 7828 21238 7840
rect 21269 7837 21281 7840
rect 21315 7868 21327 7871
rect 21634 7868 21640 7880
rect 21315 7840 21640 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 16632 7772 16896 7800
rect 16945 7803 17003 7809
rect 16632 7760 16638 7772
rect 16945 7769 16957 7803
rect 16991 7769 17003 7803
rect 16945 7763 17003 7769
rect 10836 7704 11192 7732
rect 11977 7735 12035 7741
rect 10836 7692 10842 7704
rect 11977 7701 11989 7735
rect 12023 7701 12035 7735
rect 11977 7695 12035 7701
rect 14093 7735 14151 7741
rect 14093 7701 14105 7735
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 15378 7692 15384 7744
rect 15436 7732 15442 7744
rect 16206 7732 16212 7744
rect 15436 7704 16212 7732
rect 15436 7692 15442 7704
rect 16206 7692 16212 7704
rect 16264 7732 16270 7744
rect 16960 7732 16988 7763
rect 19518 7760 19524 7812
rect 19576 7800 19582 7812
rect 19812 7800 19840 7828
rect 20438 7800 20444 7812
rect 19576 7772 20444 7800
rect 19576 7760 19582 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 21744 7800 21772 7831
rect 22186 7828 22192 7880
rect 22244 7828 22250 7880
rect 22830 7828 22836 7880
rect 22888 7868 22894 7880
rect 23385 7871 23443 7877
rect 23385 7868 23397 7871
rect 22888 7840 23397 7868
rect 22888 7828 22894 7840
rect 23385 7837 23397 7840
rect 23431 7837 23443 7871
rect 23385 7831 23443 7837
rect 24489 7871 24547 7877
rect 24489 7837 24501 7871
rect 24535 7837 24547 7871
rect 24489 7831 24547 7837
rect 20864 7772 21772 7800
rect 20864 7760 20870 7772
rect 22462 7760 22468 7812
rect 22520 7800 22526 7812
rect 22925 7803 22983 7809
rect 22925 7800 22937 7803
rect 22520 7772 22937 7800
rect 22520 7760 22526 7772
rect 22925 7769 22937 7772
rect 22971 7800 22983 7803
rect 24504 7800 24532 7831
rect 22971 7772 24532 7800
rect 22971 7769 22983 7772
rect 22925 7763 22983 7769
rect 24670 7760 24676 7812
rect 24728 7800 24734 7812
rect 24765 7803 24823 7809
rect 24765 7800 24777 7803
rect 24728 7772 24777 7800
rect 24728 7760 24734 7772
rect 24765 7769 24777 7772
rect 24811 7769 24823 7803
rect 24765 7763 24823 7769
rect 25774 7760 25780 7812
rect 25832 7760 25838 7812
rect 16264 7704 16988 7732
rect 16264 7692 16270 7704
rect 1104 7642 26864 7664
rect 1104 7590 3658 7642
rect 3710 7590 3722 7642
rect 3774 7590 3786 7642
rect 3838 7590 3850 7642
rect 3902 7590 3914 7642
rect 3966 7590 3978 7642
rect 4030 7590 7658 7642
rect 7710 7590 7722 7642
rect 7774 7590 7786 7642
rect 7838 7590 7850 7642
rect 7902 7590 7914 7642
rect 7966 7590 7978 7642
rect 8030 7590 11658 7642
rect 11710 7590 11722 7642
rect 11774 7590 11786 7642
rect 11838 7590 11850 7642
rect 11902 7590 11914 7642
rect 11966 7590 11978 7642
rect 12030 7590 15658 7642
rect 15710 7590 15722 7642
rect 15774 7590 15786 7642
rect 15838 7590 15850 7642
rect 15902 7590 15914 7642
rect 15966 7590 15978 7642
rect 16030 7590 19658 7642
rect 19710 7590 19722 7642
rect 19774 7590 19786 7642
rect 19838 7590 19850 7642
rect 19902 7590 19914 7642
rect 19966 7590 19978 7642
rect 20030 7590 23658 7642
rect 23710 7590 23722 7642
rect 23774 7590 23786 7642
rect 23838 7590 23850 7642
rect 23902 7590 23914 7642
rect 23966 7590 23978 7642
rect 24030 7590 26864 7642
rect 1104 7568 26864 7590
rect 2593 7531 2651 7537
rect 2593 7497 2605 7531
rect 2639 7528 2651 7531
rect 2774 7528 2780 7540
rect 2639 7500 2780 7528
rect 2639 7497 2651 7500
rect 2593 7491 2651 7497
rect 2774 7488 2780 7500
rect 2832 7528 2838 7540
rect 2832 7500 4200 7528
rect 2832 7488 2838 7500
rect 3421 7463 3479 7469
rect 3421 7429 3433 7463
rect 3467 7460 3479 7463
rect 3510 7460 3516 7472
rect 3467 7432 3516 7460
rect 3467 7429 3479 7432
rect 3421 7423 3479 7429
rect 3510 7420 3516 7432
rect 3568 7460 3574 7472
rect 3568 7432 3924 7460
rect 3568 7420 3574 7432
rect 3896 7401 3924 7432
rect 4062 7420 4068 7472
rect 4120 7420 4126 7472
rect 4172 7469 4200 7500
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 5445 7531 5503 7537
rect 5445 7528 5457 7531
rect 4580 7500 5457 7528
rect 4580 7488 4586 7500
rect 5445 7497 5457 7500
rect 5491 7528 5503 7531
rect 5718 7528 5724 7540
rect 5491 7500 5724 7528
rect 5491 7497 5503 7500
rect 5445 7491 5503 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 7374 7528 7380 7540
rect 7331 7500 7380 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 7653 7531 7711 7537
rect 7653 7497 7665 7531
rect 7699 7528 7711 7531
rect 8110 7528 8116 7540
rect 7699 7500 8116 7528
rect 7699 7497 7711 7500
rect 7653 7491 7711 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 9180 7500 9689 7528
rect 9180 7488 9186 7500
rect 9677 7497 9689 7500
rect 9723 7497 9735 7531
rect 9677 7491 9735 7497
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10778 7528 10784 7540
rect 10091 7500 10784 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 13173 7531 13231 7537
rect 13173 7528 13185 7531
rect 12676 7500 13185 7528
rect 12676 7488 12682 7500
rect 13173 7497 13185 7500
rect 13219 7497 13231 7531
rect 13173 7491 13231 7497
rect 13262 7488 13268 7540
rect 13320 7488 13326 7540
rect 13630 7488 13636 7540
rect 13688 7488 13694 7540
rect 13722 7488 13728 7540
rect 13780 7488 13786 7540
rect 14369 7531 14427 7537
rect 14369 7497 14381 7531
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 4157 7463 4215 7469
rect 4157 7429 4169 7463
rect 4203 7429 4215 7463
rect 4157 7423 4215 7429
rect 4264 7432 8432 7460
rect 4264 7401 4292 7432
rect 8404 7404 8432 7432
rect 10134 7420 10140 7472
rect 10192 7420 10198 7472
rect 12066 7469 12072 7472
rect 12060 7460 12072 7469
rect 12027 7432 12072 7460
rect 12060 7423 12072 7432
rect 12066 7420 12072 7423
rect 12124 7420 12130 7472
rect 14384 7460 14412 7491
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 16485 7531 16543 7537
rect 14608 7500 16436 7528
rect 14608 7488 14614 7500
rect 15350 7463 15408 7469
rect 15350 7460 15362 7463
rect 14384 7432 15362 7460
rect 15350 7429 15362 7432
rect 15396 7429 15408 7463
rect 16408 7460 16436 7500
rect 16485 7497 16497 7531
rect 16531 7528 16543 7531
rect 16758 7528 16764 7540
rect 16531 7500 16764 7528
rect 16531 7497 16543 7500
rect 16485 7491 16543 7497
rect 16758 7488 16764 7500
rect 16816 7528 16822 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16816 7500 17049 7528
rect 16816 7488 16822 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17586 7528 17592 7540
rect 17184 7500 17592 7528
rect 17184 7488 17190 7500
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 23109 7531 23167 7537
rect 19484 7500 20300 7528
rect 19484 7488 19490 7500
rect 18414 7460 18420 7472
rect 16408 7432 18420 7460
rect 15350 7423 15408 7429
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 18506 7420 18512 7472
rect 18564 7460 18570 7472
rect 19889 7463 19947 7469
rect 19889 7460 19901 7463
rect 18564 7432 19901 7460
rect 18564 7420 18570 7432
rect 19889 7429 19901 7432
rect 19935 7429 19947 7463
rect 19889 7423 19947 7429
rect 20272 7460 20300 7500
rect 21468 7500 22232 7528
rect 20272 7432 21036 7460
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3881 7395 3939 7401
rect 2731 7364 3556 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 3528 7333 3556 7364
rect 3881 7361 3893 7395
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 5442 7392 5448 7404
rect 5307 7364 5448 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7392 7067 7395
rect 7558 7392 7564 7404
rect 7055 7364 7564 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 8113 7395 8171 7401
rect 7668 7364 7880 7392
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 3513 7327 3571 7333
rect 2915 7296 3464 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 1854 7216 1860 7268
rect 1912 7256 1918 7268
rect 3053 7259 3111 7265
rect 3053 7256 3065 7259
rect 1912 7228 3065 7256
rect 1912 7216 1918 7228
rect 3053 7225 3065 7228
rect 3099 7225 3111 7259
rect 3436 7256 3464 7296
rect 3513 7293 3525 7327
rect 3559 7324 3571 7327
rect 3602 7324 3608 7336
rect 3559 7296 3608 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 4614 7324 4620 7336
rect 3743 7296 4620 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 4614 7284 4620 7296
rect 4672 7324 4678 7336
rect 6178 7324 6184 7336
rect 4672 7296 6184 7324
rect 4672 7284 4678 7296
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 7668 7324 7696 7364
rect 6880 7296 7696 7324
rect 6880 7284 6886 7296
rect 7742 7284 7748 7336
rect 7800 7284 7806 7336
rect 7852 7333 7880 7364
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 8018 7324 8024 7336
rect 7883 7296 8024 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8128 7324 8156 7355
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 8478 7352 8484 7404
rect 8536 7352 8542 7404
rect 8570 7352 8576 7404
rect 8628 7401 8634 7404
rect 8628 7355 8636 7401
rect 10594 7392 10600 7404
rect 10060 7364 10600 7392
rect 8628 7352 8634 7355
rect 10060 7324 10088 7364
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 13998 7392 14004 7404
rect 11020 7364 14004 7392
rect 11020 7352 11026 7364
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14185 7395 14243 7401
rect 14185 7361 14197 7395
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 8128 7296 10088 7324
rect 10318 7284 10324 7336
rect 10376 7284 10382 7336
rect 11514 7284 11520 7336
rect 11572 7324 11578 7336
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11572 7296 11805 7324
rect 11572 7284 11578 7296
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 13504 7296 13829 7324
rect 13504 7284 13510 7296
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 8294 7256 8300 7268
rect 3436 7228 8300 7256
rect 3053 7219 3111 7225
rect 8294 7216 8300 7228
rect 8352 7256 8358 7268
rect 11238 7256 11244 7268
rect 8352 7228 11244 7256
rect 8352 7216 8358 7228
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 2225 7191 2283 7197
rect 2225 7188 2237 7191
rect 1728 7160 2237 7188
rect 1728 7148 1734 7160
rect 2225 7157 2237 7160
rect 2271 7157 2283 7191
rect 2225 7151 2283 7157
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 5258 7188 5264 7200
rect 4479 7160 5264 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 6730 7148 6736 7200
rect 6788 7188 6794 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6788 7160 6837 7188
rect 6788 7148 6794 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 8754 7148 8760 7200
rect 8812 7148 8818 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10318 7188 10324 7200
rect 10008 7160 10324 7188
rect 10008 7148 10014 7160
rect 10318 7148 10324 7160
rect 10376 7188 10382 7200
rect 14090 7188 14096 7200
rect 10376 7160 14096 7188
rect 10376 7148 10382 7160
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 14200 7188 14228 7355
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 14884 7364 15117 7392
rect 14884 7352 14890 7364
rect 15105 7361 15117 7364
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18656 7364 18889 7392
rect 18656 7352 18662 7364
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7392 19487 7395
rect 19518 7392 19524 7404
rect 19475 7364 19524 7392
rect 19475 7361 19487 7364
rect 19429 7355 19487 7361
rect 17310 7284 17316 7336
rect 17368 7284 17374 7336
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 17828 7296 18429 7324
rect 17828 7284 17834 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 18690 7284 18696 7336
rect 18748 7324 18754 7336
rect 18984 7324 19012 7355
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 20070 7392 20076 7404
rect 19659 7364 20076 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20272 7392 20300 7432
rect 20349 7395 20407 7401
rect 20349 7392 20361 7395
rect 20272 7364 20361 7392
rect 20349 7361 20361 7364
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 20438 7352 20444 7404
rect 20496 7352 20502 7404
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7361 20959 7395
rect 21008 7392 21036 7432
rect 21266 7420 21272 7472
rect 21324 7460 21330 7472
rect 21468 7460 21496 7500
rect 21324 7432 21496 7460
rect 22204 7460 22232 7500
rect 23109 7497 23121 7531
rect 23155 7528 23167 7531
rect 25130 7528 25136 7540
rect 23155 7500 25136 7528
rect 23155 7497 23167 7500
rect 23109 7491 23167 7497
rect 25130 7488 25136 7500
rect 25188 7528 25194 7540
rect 25406 7528 25412 7540
rect 25188 7500 25412 7528
rect 25188 7488 25194 7500
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 26510 7488 26516 7540
rect 26568 7488 26574 7540
rect 22204 7432 22692 7460
rect 21324 7420 21330 7432
rect 21468 7401 21496 7432
rect 21453 7395 21511 7401
rect 21008 7364 21404 7392
rect 20901 7355 20959 7361
rect 18748 7296 19012 7324
rect 18748 7284 18754 7296
rect 19702 7284 19708 7336
rect 19760 7324 19766 7336
rect 19797 7327 19855 7333
rect 19797 7324 19809 7327
rect 19760 7296 19809 7324
rect 19760 7284 19766 7296
rect 19797 7293 19809 7296
rect 19843 7324 19855 7327
rect 20162 7324 20168 7336
rect 19843 7296 20168 7324
rect 19843 7293 19855 7296
rect 19797 7287 19855 7293
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 20714 7284 20720 7336
rect 20772 7324 20778 7336
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 20772 7296 20821 7324
rect 20772 7284 20778 7296
rect 20809 7293 20821 7296
rect 20855 7293 20867 7327
rect 20916 7324 20944 7355
rect 21082 7324 21088 7336
rect 20916 7296 21088 7324
rect 20809 7287 20867 7293
rect 21082 7284 21088 7296
rect 21140 7284 21146 7336
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7293 21327 7327
rect 21376 7324 21404 7364
rect 21453 7361 21465 7395
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 21637 7395 21695 7401
rect 21637 7361 21649 7395
rect 21683 7392 21695 7395
rect 22370 7392 22376 7404
rect 21683 7364 22376 7392
rect 21683 7361 21695 7364
rect 21637 7355 21695 7361
rect 21652 7324 21680 7355
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 22664 7401 22692 7432
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22738 7352 22744 7404
rect 22796 7352 22802 7404
rect 23477 7395 23535 7401
rect 23477 7392 23489 7395
rect 22848 7364 23489 7392
rect 21376 7296 21680 7324
rect 21269 7287 21327 7293
rect 16390 7216 16396 7268
rect 16448 7256 16454 7268
rect 20180 7256 20208 7284
rect 21284 7256 21312 7287
rect 21726 7284 21732 7336
rect 21784 7324 21790 7336
rect 22848 7324 22876 7364
rect 23477 7361 23489 7364
rect 23523 7361 23535 7395
rect 23477 7355 23535 7361
rect 23566 7352 23572 7404
rect 23624 7392 23630 7404
rect 23753 7395 23811 7401
rect 23753 7392 23765 7395
rect 23624 7364 23765 7392
rect 23624 7352 23630 7364
rect 23753 7361 23765 7364
rect 23799 7361 23811 7395
rect 23753 7355 23811 7361
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 24912 7364 25053 7392
rect 24912 7352 24918 7364
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 26326 7352 26332 7404
rect 26384 7352 26390 7404
rect 21784 7296 22876 7324
rect 22925 7327 22983 7333
rect 21784 7284 21790 7296
rect 22925 7293 22937 7327
rect 22971 7293 22983 7327
rect 22925 7287 22983 7293
rect 16448 7228 16804 7256
rect 20180 7228 21312 7256
rect 16448 7216 16454 7228
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 14200 7160 16681 7188
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16776 7188 16804 7228
rect 18782 7188 18788 7200
rect 16776 7160 18788 7188
rect 16669 7151 16727 7157
rect 18782 7148 18788 7160
rect 18840 7188 18846 7200
rect 20346 7188 20352 7200
rect 18840 7160 20352 7188
rect 18840 7148 18846 7160
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 20438 7148 20444 7200
rect 20496 7188 20502 7200
rect 20898 7188 20904 7200
rect 20496 7160 20904 7188
rect 20496 7148 20502 7160
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 21284 7188 21312 7228
rect 21634 7216 21640 7268
rect 21692 7216 21698 7268
rect 22370 7216 22376 7268
rect 22428 7256 22434 7268
rect 22738 7256 22744 7268
rect 22428 7228 22744 7256
rect 22428 7216 22434 7228
rect 22738 7216 22744 7228
rect 22796 7216 22802 7268
rect 22094 7188 22100 7200
rect 21284 7160 22100 7188
rect 22094 7148 22100 7160
rect 22152 7188 22158 7200
rect 22940 7188 22968 7287
rect 24670 7284 24676 7336
rect 24728 7284 24734 7336
rect 25130 7284 25136 7336
rect 25188 7284 25194 7336
rect 22152 7160 22968 7188
rect 22152 7148 22158 7160
rect 1104 7098 26864 7120
rect 1104 7046 2918 7098
rect 2970 7046 2982 7098
rect 3034 7046 3046 7098
rect 3098 7046 3110 7098
rect 3162 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 6918 7098
rect 6970 7046 6982 7098
rect 7034 7046 7046 7098
rect 7098 7046 7110 7098
rect 7162 7046 7174 7098
rect 7226 7046 7238 7098
rect 7290 7046 10918 7098
rect 10970 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 11238 7098
rect 11290 7046 14918 7098
rect 14970 7046 14982 7098
rect 15034 7046 15046 7098
rect 15098 7046 15110 7098
rect 15162 7046 15174 7098
rect 15226 7046 15238 7098
rect 15290 7046 18918 7098
rect 18970 7046 18982 7098
rect 19034 7046 19046 7098
rect 19098 7046 19110 7098
rect 19162 7046 19174 7098
rect 19226 7046 19238 7098
rect 19290 7046 22918 7098
rect 22970 7046 22982 7098
rect 23034 7046 23046 7098
rect 23098 7046 23110 7098
rect 23162 7046 23174 7098
rect 23226 7046 23238 7098
rect 23290 7046 26864 7098
rect 1104 7024 26864 7046
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 6822 6984 6828 6996
rect 5224 6956 6828 6984
rect 5224 6944 5230 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7616 6956 7941 6984
rect 7616 6944 7622 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 7929 6947 7987 6953
rect 8018 6944 8024 6996
rect 8076 6984 8082 6996
rect 10778 6984 10784 6996
rect 8076 6956 10784 6984
rect 8076 6944 8082 6956
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 11422 6944 11428 6996
rect 11480 6984 11486 6996
rect 14642 6984 14648 6996
rect 11480 6956 14648 6984
rect 11480 6944 11486 6956
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 15378 6984 15384 6996
rect 15028 6956 15384 6984
rect 7837 6919 7895 6925
rect 7837 6885 7849 6919
rect 7883 6916 7895 6919
rect 8202 6916 8208 6928
rect 7883 6888 8208 6916
rect 7883 6885 7895 6888
rect 7837 6879 7895 6885
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 8294 6876 8300 6928
rect 8352 6876 8358 6928
rect 8386 6876 8392 6928
rect 8444 6916 8450 6928
rect 15028 6916 15056 6956
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 16393 6987 16451 6993
rect 16393 6953 16405 6987
rect 16439 6984 16451 6987
rect 16482 6984 16488 6996
rect 16439 6956 16488 6984
rect 16439 6953 16451 6956
rect 16393 6947 16451 6953
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 18782 6944 18788 6996
rect 18840 6984 18846 6996
rect 19337 6987 19395 6993
rect 19337 6984 19349 6987
rect 18840 6956 19349 6984
rect 18840 6944 18846 6956
rect 19337 6953 19349 6956
rect 19383 6953 19395 6987
rect 19337 6947 19395 6953
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 20438 6984 20444 6996
rect 19576 6956 20444 6984
rect 19576 6944 19582 6956
rect 20438 6944 20444 6956
rect 20496 6984 20502 6996
rect 20496 6956 21864 6984
rect 20496 6944 20502 6956
rect 8444 6888 15056 6916
rect 19306 6888 20300 6916
rect 8444 6876 8450 6888
rect 8312 6848 8340 6876
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 5184 6820 6500 6848
rect 8312 6820 8493 6848
rect 1394 6740 1400 6792
rect 1452 6740 1458 6792
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1854 6780 1860 6792
rect 1719 6752 1860 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 1946 6740 1952 6792
rect 2004 6780 2010 6792
rect 2004 6752 2360 6780
rect 2004 6740 2010 6752
rect 2194 6715 2252 6721
rect 2194 6712 2206 6715
rect 1596 6684 2206 6712
rect 1596 6653 1624 6684
rect 2194 6681 2206 6684
rect 2240 6681 2252 6715
rect 2332 6712 2360 6752
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6780 3847 6783
rect 5184 6780 5212 6820
rect 6472 6792 6500 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6848 18291 6851
rect 19306 6848 19334 6888
rect 18279 6820 19334 6848
rect 20272 6848 20300 6888
rect 20898 6876 20904 6928
rect 20956 6916 20962 6928
rect 21266 6916 21272 6928
rect 20956 6888 21272 6916
rect 20956 6876 20962 6888
rect 21266 6876 21272 6888
rect 21324 6876 21330 6928
rect 20714 6848 20720 6860
rect 20272 6820 20720 6848
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 3835 6752 5212 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 3804 6712 3832 6743
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 5629 6783 5687 6789
rect 5629 6780 5641 6783
rect 5460 6752 5641 6780
rect 4034 6715 4092 6721
rect 4034 6712 4046 6715
rect 2332 6684 3832 6712
rect 3896 6684 4046 6712
rect 2194 6675 2252 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 1854 6604 1860 6656
rect 1912 6604 1918 6656
rect 3326 6604 3332 6656
rect 3384 6604 3390 6656
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3896 6644 3924 6684
rect 4034 6681 4046 6684
rect 4080 6681 4092 6715
rect 4034 6675 4092 6681
rect 3651 6616 3924 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 4764 6616 5181 6644
rect 4764 6604 4770 6616
rect 5169 6613 5181 6616
rect 5215 6644 5227 6647
rect 5460 6644 5488 6752
rect 5629 6749 5641 6752
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 5767 6783 5825 6789
rect 5767 6749 5779 6783
rect 5813 6780 5825 6783
rect 6362 6780 6368 6792
rect 5813 6752 6368 6780
rect 5813 6749 5825 6752
rect 5767 6743 5825 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 6730 6789 6736 6792
rect 6724 6780 6736 6789
rect 6691 6752 6736 6780
rect 6724 6743 6736 6752
rect 6730 6740 6736 6743
rect 6788 6740 6794 6792
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 8260 6752 8309 6780
rect 8260 6740 8266 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8662 6780 8668 6792
rect 8435 6752 8668 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9916 6752 10057 6780
rect 9916 6740 9922 6752
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 14826 6740 14832 6792
rect 14884 6780 14890 6792
rect 15013 6783 15071 6789
rect 15013 6780 15025 6783
rect 14884 6752 15025 6780
rect 14884 6740 14890 6752
rect 15013 6749 15025 6752
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 15280 6783 15338 6789
rect 15280 6749 15292 6783
rect 15326 6780 15338 6783
rect 15562 6780 15568 6792
rect 15326 6752 15568 6780
rect 15326 6749 15338 6752
rect 15280 6743 15338 6749
rect 15562 6740 15568 6752
rect 15620 6740 15626 6792
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6712 5595 6715
rect 13538 6712 13544 6724
rect 5583 6684 6316 6712
rect 5583 6681 5595 6684
rect 5537 6675 5595 6681
rect 5215 6616 5488 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5902 6604 5908 6656
rect 5960 6604 5966 6656
rect 6288 6644 6316 6684
rect 7576 6684 13544 6712
rect 7576 6644 7604 6684
rect 13538 6672 13544 6684
rect 13596 6712 13602 6724
rect 16574 6712 16580 6724
rect 13596 6684 16580 6712
rect 13596 6672 13602 6684
rect 16574 6672 16580 6684
rect 16632 6672 16638 6724
rect 6288 6616 7604 6644
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 9674 6644 9680 6656
rect 8168 6616 9680 6644
rect 8168 6604 8174 6616
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 9861 6647 9919 6653
rect 9861 6644 9873 6647
rect 9824 6616 9873 6644
rect 9824 6604 9830 6616
rect 9861 6613 9873 6616
rect 9907 6613 9919 6647
rect 18340 6644 18368 6743
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19702 6780 19708 6792
rect 19107 6752 19708 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 19794 6740 19800 6792
rect 19852 6740 19858 6792
rect 20272 6789 20300 6820
rect 20714 6808 20720 6820
rect 20772 6848 20778 6860
rect 21836 6848 21864 6956
rect 21910 6944 21916 6996
rect 21968 6984 21974 6996
rect 22465 6987 22523 6993
rect 22465 6984 22477 6987
rect 21968 6956 22477 6984
rect 21968 6944 21974 6956
rect 22465 6953 22477 6956
rect 22511 6953 22523 6987
rect 22465 6947 22523 6953
rect 25222 6944 25228 6996
rect 25280 6944 25286 6996
rect 24673 6851 24731 6857
rect 20772 6820 21772 6848
rect 21836 6820 22232 6848
rect 20772 6808 20778 6820
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 20441 6783 20499 6789
rect 20441 6749 20453 6783
rect 20487 6780 20499 6783
rect 20530 6780 20536 6792
rect 20487 6752 20536 6780
rect 20487 6749 20499 6752
rect 20441 6743 20499 6749
rect 18693 6715 18751 6721
rect 18693 6681 18705 6715
rect 18739 6712 18751 6715
rect 19242 6712 19248 6724
rect 18739 6684 19248 6712
rect 18739 6681 18751 6684
rect 18693 6675 18751 6681
rect 19242 6672 19248 6684
rect 19300 6672 19306 6724
rect 19426 6672 19432 6724
rect 19484 6712 19490 6724
rect 19996 6712 20024 6743
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20622 6740 20628 6792
rect 20680 6740 20686 6792
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21192 6712 21220 6743
rect 21266 6740 21272 6792
rect 21324 6740 21330 6792
rect 21634 6740 21640 6792
rect 21692 6740 21698 6792
rect 21744 6789 21772 6820
rect 21729 6783 21787 6789
rect 21729 6749 21741 6783
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 22094 6740 22100 6792
rect 22152 6740 22158 6792
rect 22204 6789 22232 6820
rect 24673 6817 24685 6851
rect 24719 6817 24731 6851
rect 24673 6811 24731 6817
rect 22189 6783 22247 6789
rect 22189 6749 22201 6783
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22554 6740 22560 6792
rect 22612 6780 22618 6792
rect 23106 6780 23112 6792
rect 22612 6752 23112 6780
rect 22612 6740 22618 6752
rect 23106 6740 23112 6752
rect 23164 6780 23170 6792
rect 23566 6780 23572 6792
rect 23164 6752 23572 6780
rect 23164 6740 23170 6752
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 24210 6740 24216 6792
rect 24268 6780 24274 6792
rect 24578 6780 24584 6792
rect 24268 6752 24584 6780
rect 24268 6740 24274 6752
rect 24578 6740 24584 6752
rect 24636 6740 24642 6792
rect 24688 6780 24716 6811
rect 24946 6808 24952 6860
rect 25004 6808 25010 6860
rect 25682 6808 25688 6860
rect 25740 6808 25746 6860
rect 25041 6783 25099 6789
rect 25041 6780 25053 6783
rect 24688 6752 25053 6780
rect 25041 6749 25053 6752
rect 25087 6749 25099 6783
rect 25041 6743 25099 6749
rect 25225 6783 25283 6789
rect 25225 6749 25237 6783
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 19484 6684 21220 6712
rect 19484 6672 19490 6684
rect 19334 6644 19340 6656
rect 18340 6616 19340 6644
rect 9861 6607 9919 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 20990 6604 20996 6656
rect 21048 6604 21054 6656
rect 21192 6644 21220 6684
rect 21542 6672 21548 6724
rect 21600 6712 21606 6724
rect 22456 6715 22514 6721
rect 22456 6712 22468 6715
rect 21600 6684 22468 6712
rect 21600 6672 21606 6684
rect 22456 6681 22468 6684
rect 22502 6712 22514 6715
rect 22572 6712 22600 6740
rect 22502 6684 22600 6712
rect 22502 6681 22514 6684
rect 22456 6675 22514 6681
rect 22830 6672 22836 6724
rect 22888 6672 22894 6724
rect 22186 6644 22192 6656
rect 21192 6616 22192 6644
rect 22186 6604 22192 6616
rect 22244 6644 22250 6656
rect 22554 6644 22560 6656
rect 22244 6616 22560 6644
rect 22244 6604 22250 6616
rect 22554 6604 22560 6616
rect 22612 6604 22618 6656
rect 25056 6644 25084 6743
rect 25240 6712 25268 6743
rect 25314 6740 25320 6792
rect 25372 6780 25378 6792
rect 25501 6783 25559 6789
rect 25501 6780 25513 6783
rect 25372 6752 25513 6780
rect 25372 6740 25378 6752
rect 25501 6749 25513 6752
rect 25547 6780 25559 6783
rect 25593 6783 25651 6789
rect 25593 6780 25605 6783
rect 25547 6752 25605 6780
rect 25547 6749 25559 6752
rect 25501 6743 25559 6749
rect 25593 6749 25605 6752
rect 25639 6749 25651 6783
rect 25777 6783 25835 6789
rect 25777 6780 25789 6783
rect 25593 6743 25651 6749
rect 25700 6752 25789 6780
rect 25700 6724 25728 6752
rect 25777 6749 25789 6752
rect 25823 6749 25835 6783
rect 25777 6743 25835 6749
rect 25240 6684 25636 6712
rect 25608 6656 25636 6684
rect 25682 6672 25688 6724
rect 25740 6672 25746 6724
rect 25498 6644 25504 6656
rect 25056 6616 25504 6644
rect 25498 6604 25504 6616
rect 25556 6604 25562 6656
rect 25590 6604 25596 6656
rect 25648 6604 25654 6656
rect 1104 6554 26864 6576
rect 1104 6502 3658 6554
rect 3710 6502 3722 6554
rect 3774 6502 3786 6554
rect 3838 6502 3850 6554
rect 3902 6502 3914 6554
rect 3966 6502 3978 6554
rect 4030 6502 7658 6554
rect 7710 6502 7722 6554
rect 7774 6502 7786 6554
rect 7838 6502 7850 6554
rect 7902 6502 7914 6554
rect 7966 6502 7978 6554
rect 8030 6502 11658 6554
rect 11710 6502 11722 6554
rect 11774 6502 11786 6554
rect 11838 6502 11850 6554
rect 11902 6502 11914 6554
rect 11966 6502 11978 6554
rect 12030 6502 15658 6554
rect 15710 6502 15722 6554
rect 15774 6502 15786 6554
rect 15838 6502 15850 6554
rect 15902 6502 15914 6554
rect 15966 6502 15978 6554
rect 16030 6502 19658 6554
rect 19710 6502 19722 6554
rect 19774 6502 19786 6554
rect 19838 6502 19850 6554
rect 19902 6502 19914 6554
rect 19966 6502 19978 6554
rect 20030 6502 23658 6554
rect 23710 6502 23722 6554
rect 23774 6502 23786 6554
rect 23838 6502 23850 6554
rect 23902 6502 23914 6554
rect 23966 6502 23978 6554
rect 24030 6502 26864 6554
rect 1104 6480 26864 6502
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 3476 6412 4353 6440
rect 3476 6400 3482 6412
rect 4341 6409 4353 6412
rect 4387 6409 4399 6443
rect 4341 6403 4399 6409
rect 4706 6400 4712 6452
rect 4764 6400 4770 6452
rect 4801 6443 4859 6449
rect 4801 6409 4813 6443
rect 4847 6440 4859 6443
rect 5442 6440 5448 6452
rect 4847 6412 5448 6440
rect 4847 6409 4859 6412
rect 4801 6403 4859 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 7745 6443 7803 6449
rect 7745 6409 7757 6443
rect 7791 6440 7803 6443
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 7791 6412 8217 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 8205 6409 8217 6412
rect 8251 6440 8263 6443
rect 8478 6440 8484 6452
rect 8251 6412 8484 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 9398 6400 9404 6452
rect 9456 6400 9462 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10284 6412 10885 6440
rect 10284 6400 10290 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 12897 6443 12955 6449
rect 12897 6409 12909 6443
rect 12943 6440 12955 6443
rect 13354 6440 13360 6452
rect 12943 6412 13360 6440
rect 12943 6409 12955 6412
rect 12897 6403 12955 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 13722 6440 13728 6452
rect 13495 6412 13728 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 16206 6400 16212 6452
rect 16264 6440 16270 6452
rect 18782 6440 18788 6452
rect 16264 6412 18788 6440
rect 16264 6400 16270 6412
rect 18782 6400 18788 6412
rect 18840 6400 18846 6452
rect 19981 6443 20039 6449
rect 19981 6409 19993 6443
rect 20027 6440 20039 6443
rect 20162 6440 20168 6452
rect 20027 6412 20168 6440
rect 20027 6409 20039 6412
rect 19981 6403 20039 6409
rect 20162 6400 20168 6412
rect 20220 6400 20226 6452
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20312 6412 21189 6440
rect 20312 6400 20318 6412
rect 21177 6409 21189 6412
rect 21223 6440 21235 6443
rect 21634 6440 21640 6452
rect 21223 6412 21640 6440
rect 21223 6409 21235 6412
rect 21177 6403 21235 6409
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 21726 6400 21732 6452
rect 21784 6440 21790 6452
rect 22649 6443 22707 6449
rect 22649 6440 22661 6443
rect 21784 6412 22661 6440
rect 21784 6400 21790 6412
rect 22649 6409 22661 6412
rect 22695 6409 22707 6443
rect 22649 6403 22707 6409
rect 23293 6443 23351 6449
rect 23293 6409 23305 6443
rect 23339 6440 23351 6443
rect 23382 6440 23388 6452
rect 23339 6412 23388 6440
rect 23339 6409 23351 6412
rect 23293 6403 23351 6409
rect 1854 6332 1860 6384
rect 1912 6372 1918 6384
rect 2194 6375 2252 6381
rect 2194 6372 2206 6375
rect 1912 6344 2206 6372
rect 1912 6332 1918 6344
rect 2194 6341 2206 6344
rect 2240 6341 2252 6375
rect 2194 6335 2252 6341
rect 3326 6332 3332 6384
rect 3384 6372 3390 6384
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3384 6344 3801 6372
rect 3384 6332 3390 6344
rect 3789 6341 3801 6344
rect 3835 6372 3847 6375
rect 5350 6372 5356 6384
rect 3835 6344 5356 6372
rect 3835 6341 3847 6344
rect 3789 6335 3847 6341
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 6454 6372 6460 6384
rect 6380 6344 6460 6372
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 1946 6264 1952 6316
rect 2004 6264 2010 6316
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 4522 6304 4528 6316
rect 3927 6276 4528 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 6380 6313 6408 6344
rect 6454 6332 6460 6344
rect 6512 6372 6518 6384
rect 6822 6372 6828 6384
rect 6512 6344 6828 6372
rect 6512 6332 6518 6344
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 8297 6375 8355 6381
rect 8297 6341 8309 6375
rect 8343 6372 8355 6375
rect 8662 6372 8668 6384
rect 8343 6344 8668 6372
rect 8343 6341 8355 6344
rect 8297 6335 8355 6341
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 8941 6375 8999 6381
rect 8941 6372 8953 6375
rect 8812 6344 8953 6372
rect 8812 6332 8818 6344
rect 8941 6341 8953 6344
rect 8987 6341 8999 6375
rect 8941 6335 8999 6341
rect 9508 6344 11284 6372
rect 9508 6316 9536 6344
rect 6638 6313 6644 6316
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6632 6267 6644 6313
rect 6638 6264 6644 6267
rect 6696 6264 6702 6316
rect 9214 6264 9220 6316
rect 9272 6264 9278 6316
rect 9490 6264 9496 6316
rect 9548 6264 9554 6316
rect 9766 6313 9772 6316
rect 9760 6304 9772 6313
rect 9727 6276 9772 6304
rect 9760 6267 9772 6276
rect 9766 6264 9772 6267
rect 9824 6264 9830 6316
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6205 5043 6239
rect 4985 6199 5043 6205
rect 1394 6128 1400 6180
rect 1452 6168 1458 6180
rect 3421 6171 3479 6177
rect 3421 6168 3433 6171
rect 1452 6140 1992 6168
rect 1452 6128 1458 6140
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1820 6072 1869 6100
rect 1820 6060 1826 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 1964 6100 1992 6140
rect 3068 6140 3433 6168
rect 3068 6100 3096 6140
rect 3421 6137 3433 6140
rect 3467 6137 3479 6171
rect 3421 6131 3479 6137
rect 1964 6072 3096 6100
rect 3329 6103 3387 6109
rect 1857 6063 1915 6069
rect 3329 6069 3341 6103
rect 3375 6100 3387 6103
rect 3510 6100 3516 6112
rect 3375 6072 3516 6100
rect 3375 6069 3387 6072
rect 3329 6063 3387 6069
rect 3510 6060 3516 6072
rect 3568 6060 3574 6112
rect 5000 6100 5028 6199
rect 7374 6196 7380 6248
rect 7432 6236 7438 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 7432 6208 8493 6236
rect 7432 6196 7438 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 8496 6168 8524 6199
rect 9030 6196 9036 6248
rect 9088 6196 9094 6248
rect 11256 6236 11284 6344
rect 17770 6332 17776 6384
rect 17828 6372 17834 6384
rect 18233 6375 18291 6381
rect 18233 6372 18245 6375
rect 17828 6344 18245 6372
rect 17828 6332 17834 6344
rect 18233 6341 18245 6344
rect 18279 6341 18291 6375
rect 20530 6372 20536 6384
rect 18233 6335 18291 6341
rect 19260 6344 20536 6372
rect 11790 6313 11796 6316
rect 11784 6267 11796 6313
rect 11790 6264 11796 6267
rect 11848 6264 11854 6316
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18656 6276 18705 6304
rect 18656 6264 18662 6276
rect 18693 6273 18705 6276
rect 18739 6273 18751 6307
rect 18693 6267 18751 6273
rect 18782 6264 18788 6316
rect 18840 6264 18846 6316
rect 19260 6313 19288 6344
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 20622 6332 20628 6384
rect 20680 6372 20686 6384
rect 21345 6375 21403 6381
rect 20680 6344 21128 6372
rect 20680 6332 20686 6344
rect 19245 6307 19303 6313
rect 19245 6273 19257 6307
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 20165 6307 20223 6313
rect 20165 6304 20177 6307
rect 19484 6276 20177 6304
rect 19484 6264 19490 6276
rect 20165 6273 20177 6276
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 20303 6276 20392 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 11514 6236 11520 6248
rect 11256 6208 11520 6236
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13596 6208 13645 6236
rect 13596 6196 13602 6208
rect 13633 6205 13645 6208
rect 13679 6236 13691 6239
rect 16390 6236 16396 6248
rect 13679 6208 16396 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 19153 6239 19211 6245
rect 19153 6205 19165 6239
rect 19199 6205 19211 6239
rect 19153 6199 19211 6205
rect 19613 6239 19671 6245
rect 19613 6205 19625 6239
rect 19659 6205 19671 6239
rect 19613 6199 19671 6205
rect 8496 6140 9076 6168
rect 7558 6100 7564 6112
rect 5000 6072 7564 6100
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7834 6060 7840 6112
rect 7892 6060 7898 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8904 6072 8953 6100
rect 8904 6060 8910 6072
rect 8941 6069 8953 6072
rect 8987 6069 8999 6103
rect 9048 6100 9076 6140
rect 12912 6140 18736 6168
rect 12912 6100 12940 6140
rect 9048 6072 12940 6100
rect 8941 6063 8999 6069
rect 12986 6060 12992 6112
rect 13044 6060 13050 6112
rect 18708 6100 18736 6140
rect 18782 6128 18788 6180
rect 18840 6168 18846 6180
rect 19168 6168 19196 6199
rect 18840 6140 19196 6168
rect 18840 6128 18846 6140
rect 19242 6128 19248 6180
rect 19300 6168 19306 6180
rect 19628 6168 19656 6199
rect 19300 6140 19656 6168
rect 20364 6168 20392 6276
rect 20714 6264 20720 6316
rect 20772 6264 20778 6316
rect 20438 6196 20444 6248
rect 20496 6236 20502 6248
rect 21100 6245 21128 6344
rect 21345 6341 21357 6375
rect 21391 6372 21403 6375
rect 21391 6344 21496 6372
rect 21391 6341 21403 6344
rect 21345 6335 21403 6341
rect 21468 6304 21496 6344
rect 21542 6332 21548 6384
rect 21600 6332 21606 6384
rect 23308 6372 23336 6403
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 23566 6400 23572 6452
rect 23624 6400 23630 6452
rect 24854 6440 24860 6452
rect 24136 6412 24860 6440
rect 22480 6344 23336 6372
rect 23477 6375 23535 6381
rect 21910 6304 21916 6316
rect 21468 6276 21916 6304
rect 21910 6264 21916 6276
rect 21968 6264 21974 6316
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 22278 6264 22284 6316
rect 22336 6264 22342 6316
rect 22480 6313 22508 6344
rect 23477 6341 23489 6375
rect 23523 6372 23535 6375
rect 24136 6372 24164 6412
rect 24854 6400 24860 6412
rect 24912 6440 24918 6452
rect 25406 6440 25412 6452
rect 25464 6449 25470 6452
rect 25464 6443 25483 6449
rect 24912 6412 25412 6440
rect 24912 6400 24918 6412
rect 25406 6400 25412 6412
rect 25471 6409 25483 6443
rect 25869 6443 25927 6449
rect 25869 6440 25881 6443
rect 25464 6403 25483 6409
rect 25516 6412 25881 6440
rect 25464 6400 25470 6403
rect 23523 6344 24164 6372
rect 23523 6341 23535 6344
rect 23477 6335 23535 6341
rect 22465 6307 22523 6313
rect 22465 6273 22477 6307
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 22830 6264 22836 6316
rect 22888 6264 22894 6316
rect 23106 6264 23112 6316
rect 23164 6264 23170 6316
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 20496 6208 20637 6236
rect 20496 6196 20502 6208
rect 20625 6205 20637 6208
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 21085 6239 21143 6245
rect 21085 6205 21097 6239
rect 21131 6236 21143 6239
rect 22296 6236 22324 6264
rect 21131 6208 22324 6236
rect 21131 6205 21143 6208
rect 21085 6199 21143 6205
rect 22646 6196 22652 6248
rect 22704 6236 22710 6248
rect 22741 6239 22799 6245
rect 22741 6236 22753 6239
rect 22704 6208 22753 6236
rect 22704 6196 22710 6208
rect 22741 6205 22753 6208
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 22848 6236 22876 6264
rect 23492 6236 23520 6335
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6304 23719 6307
rect 23845 6307 23903 6313
rect 23707 6276 23796 6304
rect 23707 6273 23719 6276
rect 23661 6267 23719 6273
rect 22848 6208 23520 6236
rect 20898 6168 20904 6180
rect 20364 6140 20904 6168
rect 19300 6128 19306 6140
rect 19628 6112 19656 6140
rect 20898 6128 20904 6140
rect 20956 6128 20962 6180
rect 22848 6168 22876 6208
rect 21376 6140 22876 6168
rect 21376 6112 21404 6140
rect 19150 6100 19156 6112
rect 18708 6072 19156 6100
rect 19150 6060 19156 6072
rect 19208 6100 19214 6112
rect 19426 6100 19432 6112
rect 19208 6072 19432 6100
rect 19208 6060 19214 6072
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 20806 6100 20812 6112
rect 19668 6072 20812 6100
rect 19668 6060 19674 6072
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 21358 6060 21364 6112
rect 21416 6060 21422 6112
rect 21821 6103 21879 6109
rect 21821 6069 21833 6103
rect 21867 6100 21879 6103
rect 21910 6100 21916 6112
rect 21867 6072 21916 6100
rect 21867 6069 21879 6072
rect 21821 6063 21879 6069
rect 21910 6060 21916 6072
rect 21968 6060 21974 6112
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 23768 6100 23796 6276
rect 23845 6273 23857 6307
rect 23891 6304 23903 6307
rect 24026 6304 24032 6316
rect 23891 6276 24032 6304
rect 23891 6273 23903 6276
rect 23845 6267 23903 6273
rect 24026 6264 24032 6276
rect 24084 6264 24090 6316
rect 24136 6313 24164 6344
rect 24302 6332 24308 6384
rect 24360 6332 24366 6384
rect 25222 6372 25228 6384
rect 24688 6344 25228 6372
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6273 24179 6307
rect 24121 6267 24179 6273
rect 24213 6307 24271 6313
rect 24213 6273 24225 6307
rect 24259 6304 24271 6307
rect 24320 6304 24348 6332
rect 24259 6276 24348 6304
rect 24397 6307 24455 6313
rect 24259 6273 24271 6276
rect 24213 6267 24271 6273
rect 24397 6273 24409 6307
rect 24443 6304 24455 6307
rect 24578 6304 24584 6316
rect 24443 6276 24584 6304
rect 24443 6273 24455 6276
rect 24397 6267 24455 6273
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 23934 6196 23940 6248
rect 23992 6196 23998 6248
rect 24305 6239 24363 6245
rect 24305 6205 24317 6239
rect 24351 6236 24363 6239
rect 24688 6236 24716 6344
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 25516 6372 25544 6412
rect 25869 6409 25881 6412
rect 25915 6409 25927 6443
rect 25869 6403 25927 6409
rect 25424 6344 25544 6372
rect 24762 6264 24768 6316
rect 24820 6264 24826 6316
rect 24351 6208 24716 6236
rect 24351 6205 24363 6208
rect 24305 6199 24363 6205
rect 24320 6100 24348 6199
rect 24854 6196 24860 6248
rect 24912 6196 24918 6248
rect 24762 6128 24768 6180
rect 24820 6168 24826 6180
rect 25424 6168 25452 6344
rect 25590 6332 25596 6384
rect 25648 6372 25654 6384
rect 25648 6344 26096 6372
rect 25648 6332 25654 6344
rect 25682 6264 25688 6316
rect 25740 6264 25746 6316
rect 25958 6264 25964 6316
rect 26016 6264 26022 6316
rect 26068 6313 26096 6344
rect 26053 6307 26111 6313
rect 26053 6273 26065 6307
rect 26099 6273 26111 6307
rect 26053 6267 26111 6273
rect 26237 6307 26295 6313
rect 26237 6273 26249 6307
rect 26283 6273 26295 6307
rect 26237 6267 26295 6273
rect 26252 6236 26280 6267
rect 25700 6208 26280 6236
rect 24820 6140 25452 6168
rect 24820 6128 24826 6140
rect 22152 6072 24348 6100
rect 22152 6060 22158 6072
rect 24854 6060 24860 6112
rect 24912 6100 24918 6112
rect 25133 6103 25191 6109
rect 25133 6100 25145 6103
rect 24912 6072 25145 6100
rect 24912 6060 24918 6072
rect 25133 6069 25145 6072
rect 25179 6100 25191 6103
rect 25314 6100 25320 6112
rect 25179 6072 25320 6100
rect 25179 6069 25191 6072
rect 25133 6063 25191 6069
rect 25314 6060 25320 6072
rect 25372 6060 25378 6112
rect 25424 6109 25452 6140
rect 25498 6128 25504 6180
rect 25556 6168 25562 6180
rect 25700 6177 25728 6208
rect 25685 6171 25743 6177
rect 25685 6168 25697 6171
rect 25556 6140 25697 6168
rect 25556 6128 25562 6140
rect 25685 6137 25697 6140
rect 25731 6137 25743 6171
rect 25685 6131 25743 6137
rect 25409 6103 25467 6109
rect 25409 6069 25421 6103
rect 25455 6069 25467 6103
rect 25409 6063 25467 6069
rect 25590 6060 25596 6112
rect 25648 6060 25654 6112
rect 26050 6060 26056 6112
rect 26108 6060 26114 6112
rect 1104 6010 26864 6032
rect 1104 5958 2918 6010
rect 2970 5958 2982 6010
rect 3034 5958 3046 6010
rect 3098 5958 3110 6010
rect 3162 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 6918 6010
rect 6970 5958 6982 6010
rect 7034 5958 7046 6010
rect 7098 5958 7110 6010
rect 7162 5958 7174 6010
rect 7226 5958 7238 6010
rect 7290 5958 10918 6010
rect 10970 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 11238 6010
rect 11290 5958 14918 6010
rect 14970 5958 14982 6010
rect 15034 5958 15046 6010
rect 15098 5958 15110 6010
rect 15162 5958 15174 6010
rect 15226 5958 15238 6010
rect 15290 5958 18918 6010
rect 18970 5958 18982 6010
rect 19034 5958 19046 6010
rect 19098 5958 19110 6010
rect 19162 5958 19174 6010
rect 19226 5958 19238 6010
rect 19290 5958 22918 6010
rect 22970 5958 22982 6010
rect 23034 5958 23046 6010
rect 23098 5958 23110 6010
rect 23162 5958 23174 6010
rect 23226 5958 23238 6010
rect 23290 5958 26864 6010
rect 1104 5936 26864 5958
rect 1946 5896 1952 5908
rect 1688 5868 1952 5896
rect 1688 5769 1716 5868
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 2832 5868 3065 5896
rect 2832 5856 2838 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 3053 5859 3111 5865
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 6733 5899 6791 5905
rect 6733 5896 6745 5899
rect 6696 5868 6745 5896
rect 6696 5856 6702 5868
rect 6733 5865 6745 5868
rect 6779 5865 6791 5899
rect 6733 5859 6791 5865
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 8662 5896 8668 5908
rect 8260 5868 8668 5896
rect 8260 5856 8266 5868
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 9858 5856 9864 5908
rect 9916 5856 9922 5908
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11848 5868 11897 5896
rect 11848 5856 11854 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 13170 5896 13176 5908
rect 11885 5859 11943 5865
rect 12406 5868 13176 5896
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 12406 5828 12434 5868
rect 13170 5856 13176 5868
rect 13228 5896 13234 5908
rect 16206 5896 16212 5908
rect 13228 5868 16212 5896
rect 13228 5856 13234 5868
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 19337 5899 19395 5905
rect 19337 5865 19349 5899
rect 19383 5896 19395 5899
rect 19426 5896 19432 5908
rect 19383 5868 19432 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 23566 5856 23572 5908
rect 23624 5896 23630 5908
rect 24029 5899 24087 5905
rect 24029 5896 24041 5899
rect 23624 5868 24041 5896
rect 23624 5856 23630 5868
rect 24029 5865 24041 5868
rect 24075 5896 24087 5899
rect 24762 5896 24768 5908
rect 24075 5868 24768 5896
rect 24075 5865 24087 5868
rect 24029 5859 24087 5865
rect 24762 5856 24768 5868
rect 24820 5856 24826 5908
rect 4120 5800 12434 5828
rect 4120 5788 4126 5800
rect 12710 5788 12716 5840
rect 12768 5828 12774 5840
rect 13449 5831 13507 5837
rect 13449 5828 13461 5831
rect 12768 5800 13461 5828
rect 12768 5788 12774 5800
rect 13449 5797 13461 5800
rect 13495 5797 13507 5831
rect 13449 5791 13507 5797
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5760 10563 5763
rect 10686 5760 10692 5772
rect 10551 5732 10692 5760
rect 10551 5729 10563 5732
rect 10505 5723 10563 5729
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 13464 5760 13492 5791
rect 16850 5788 16856 5840
rect 16908 5828 16914 5840
rect 17773 5831 17831 5837
rect 17773 5828 17785 5831
rect 16908 5800 17785 5828
rect 16908 5788 16914 5800
rect 17773 5797 17785 5800
rect 17819 5797 17831 5831
rect 18690 5828 18696 5840
rect 17773 5791 17831 5797
rect 18248 5800 18696 5828
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 13464 5732 14565 5760
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 1929 5695 1987 5701
rect 1929 5692 1941 5695
rect 1820 5664 1941 5692
rect 1820 5652 1826 5664
rect 1929 5661 1941 5664
rect 1975 5661 1987 5695
rect 1929 5655 1987 5661
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 7834 5692 7840 5704
rect 6963 5664 7840 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5692 12127 5695
rect 12986 5692 12992 5704
rect 12115 5664 12992 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5692 13691 5695
rect 13722 5692 13728 5704
rect 13679 5664 13728 5692
rect 13679 5661 13691 5664
rect 13633 5655 13691 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 13998 5652 14004 5704
rect 14056 5692 14062 5704
rect 14752 5692 14780 5723
rect 16206 5720 16212 5772
rect 16264 5720 16270 5772
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 17126 5760 17132 5772
rect 16347 5732 17132 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 18046 5692 18052 5704
rect 14056 5664 18052 5692
rect 14056 5652 14062 5664
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18248 5701 18276 5800
rect 18690 5788 18696 5800
rect 18748 5828 18754 5840
rect 20346 5828 20352 5840
rect 18748 5800 20352 5828
rect 18748 5788 18754 5800
rect 19518 5760 19524 5772
rect 18708 5732 19524 5760
rect 18708 5701 18736 5732
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 13538 5624 13544 5636
rect 7616 5596 13544 5624
rect 7616 5584 7622 5596
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 16666 5584 16672 5636
rect 16724 5624 16730 5636
rect 18432 5624 18460 5655
rect 18782 5652 18788 5704
rect 18840 5692 18846 5704
rect 18877 5695 18935 5701
rect 18877 5692 18889 5695
rect 18840 5664 18889 5692
rect 18840 5652 18846 5664
rect 18877 5661 18889 5664
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5692 19119 5695
rect 19610 5692 19616 5704
rect 19107 5664 19616 5692
rect 19107 5661 19119 5664
rect 19061 5655 19119 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 19812 5701 19840 5800
rect 20346 5788 20352 5800
rect 20404 5828 20410 5840
rect 21174 5828 21180 5840
rect 20404 5800 21180 5828
rect 20404 5788 20410 5800
rect 21174 5788 21180 5800
rect 21232 5788 21238 5840
rect 25590 5828 25596 5840
rect 22848 5800 25596 5828
rect 20625 5763 20683 5769
rect 20625 5729 20637 5763
rect 20671 5760 20683 5763
rect 20717 5763 20775 5769
rect 20717 5760 20729 5763
rect 20671 5732 20729 5760
rect 20671 5729 20683 5732
rect 20625 5723 20683 5729
rect 20717 5729 20729 5732
rect 20763 5760 20775 5763
rect 20806 5760 20812 5772
rect 20763 5732 20812 5760
rect 20763 5729 20775 5732
rect 20717 5723 20775 5729
rect 20806 5720 20812 5732
rect 20864 5720 20870 5772
rect 21726 5760 21732 5772
rect 21100 5732 21732 5760
rect 21100 5704 21128 5732
rect 21726 5720 21732 5732
rect 21784 5720 21790 5772
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 22336 5732 22692 5760
rect 22336 5720 22342 5732
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 18598 5624 18604 5636
rect 16724 5596 16988 5624
rect 18432 5596 18604 5624
rect 16724 5584 16730 5596
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 8110 5556 8116 5568
rect 6420 5528 8116 5556
rect 6420 5516 6426 5528
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 10321 5559 10379 5565
rect 10321 5556 10333 5559
rect 9456 5528 10333 5556
rect 9456 5516 9462 5528
rect 10321 5525 10333 5528
rect 10367 5525 10379 5559
rect 10321 5519 10379 5525
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 14458 5516 14464 5568
rect 14516 5516 14522 5568
rect 16390 5516 16396 5568
rect 16448 5516 16454 5568
rect 16761 5559 16819 5565
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 16850 5556 16856 5568
rect 16807 5528 16856 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 16960 5556 16988 5596
rect 18598 5584 18604 5596
rect 18656 5624 18662 5636
rect 18966 5624 18972 5636
rect 18656 5596 18972 5624
rect 18656 5584 18662 5596
rect 18966 5584 18972 5596
rect 19024 5624 19030 5636
rect 19996 5624 20024 5655
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20165 5695 20223 5701
rect 20165 5692 20177 5695
rect 20128 5664 20177 5692
rect 20128 5652 20134 5664
rect 20165 5661 20177 5664
rect 20211 5661 20223 5695
rect 20165 5655 20223 5661
rect 20254 5652 20260 5704
rect 20312 5652 20318 5704
rect 20901 5695 20959 5701
rect 20901 5661 20913 5695
rect 20947 5692 20959 5695
rect 20990 5692 20996 5704
rect 20947 5664 20996 5692
rect 20947 5661 20959 5664
rect 20901 5655 20959 5661
rect 20990 5652 20996 5664
rect 21048 5652 21054 5704
rect 21082 5652 21088 5704
rect 21140 5652 21146 5704
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 21545 5695 21603 5701
rect 21545 5692 21557 5695
rect 21232 5664 21557 5692
rect 21232 5652 21238 5664
rect 21545 5661 21557 5664
rect 21591 5661 21603 5695
rect 21545 5655 21603 5661
rect 21637 5695 21695 5701
rect 21637 5661 21649 5695
rect 21683 5692 21695 5695
rect 21818 5692 21824 5704
rect 21683 5664 21824 5692
rect 21683 5661 21695 5664
rect 21637 5655 21695 5661
rect 20438 5624 20444 5636
rect 19024 5596 20444 5624
rect 19024 5584 19030 5596
rect 20438 5584 20444 5596
rect 20496 5624 20502 5636
rect 21652 5624 21680 5655
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 22186 5652 22192 5704
rect 22244 5692 22250 5704
rect 22465 5695 22523 5701
rect 22465 5692 22477 5695
rect 22244 5664 22477 5692
rect 22244 5652 22250 5664
rect 22465 5661 22477 5664
rect 22511 5661 22523 5695
rect 22465 5655 22523 5661
rect 22554 5652 22560 5704
rect 22612 5652 22618 5704
rect 22664 5701 22692 5732
rect 22848 5701 22876 5800
rect 25590 5788 25596 5800
rect 25648 5788 25654 5840
rect 26050 5828 26056 5840
rect 25700 5800 26056 5828
rect 24854 5720 24860 5772
rect 24912 5720 24918 5772
rect 25041 5763 25099 5769
rect 25041 5729 25053 5763
rect 25087 5760 25099 5763
rect 25130 5760 25136 5772
rect 25087 5732 25136 5760
rect 25087 5729 25099 5732
rect 25041 5723 25099 5729
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 25700 5769 25728 5800
rect 26050 5788 26056 5800
rect 26108 5788 26114 5840
rect 25685 5763 25743 5769
rect 25685 5729 25697 5763
rect 25731 5729 25743 5763
rect 25685 5723 25743 5729
rect 25777 5763 25835 5769
rect 25777 5729 25789 5763
rect 25823 5729 25835 5763
rect 25777 5723 25835 5729
rect 22649 5695 22707 5701
rect 22649 5661 22661 5695
rect 22695 5661 22707 5695
rect 22649 5655 22707 5661
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5692 24271 5695
rect 24302 5692 24308 5704
rect 24259 5664 24308 5692
rect 24259 5661 24271 5664
rect 24213 5655 24271 5661
rect 24302 5652 24308 5664
rect 24360 5652 24366 5704
rect 24762 5652 24768 5704
rect 24820 5652 24826 5704
rect 20496 5596 21680 5624
rect 25148 5624 25176 5720
rect 25222 5652 25228 5704
rect 25280 5692 25286 5704
rect 25590 5692 25596 5704
rect 25280 5664 25596 5692
rect 25280 5652 25286 5664
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 25792 5624 25820 5723
rect 25148 5596 25820 5624
rect 20496 5584 20502 5596
rect 21821 5559 21879 5565
rect 21821 5556 21833 5559
rect 16960 5528 21833 5556
rect 21821 5525 21833 5528
rect 21867 5525 21879 5559
rect 21821 5519 21879 5525
rect 22186 5516 22192 5568
rect 22244 5516 22250 5568
rect 24394 5516 24400 5568
rect 24452 5516 24458 5568
rect 25222 5516 25228 5568
rect 25280 5516 25286 5568
rect 1104 5466 26864 5488
rect 1104 5414 3658 5466
rect 3710 5414 3722 5466
rect 3774 5414 3786 5466
rect 3838 5414 3850 5466
rect 3902 5414 3914 5466
rect 3966 5414 3978 5466
rect 4030 5414 7658 5466
rect 7710 5414 7722 5466
rect 7774 5414 7786 5466
rect 7838 5414 7850 5466
rect 7902 5414 7914 5466
rect 7966 5414 7978 5466
rect 8030 5414 11658 5466
rect 11710 5414 11722 5466
rect 11774 5414 11786 5466
rect 11838 5414 11850 5466
rect 11902 5414 11914 5466
rect 11966 5414 11978 5466
rect 12030 5414 15658 5466
rect 15710 5414 15722 5466
rect 15774 5414 15786 5466
rect 15838 5414 15850 5466
rect 15902 5414 15914 5466
rect 15966 5414 15978 5466
rect 16030 5414 19658 5466
rect 19710 5414 19722 5466
rect 19774 5414 19786 5466
rect 19838 5414 19850 5466
rect 19902 5414 19914 5466
rect 19966 5414 19978 5466
rect 20030 5414 23658 5466
rect 23710 5414 23722 5466
rect 23774 5414 23786 5466
rect 23838 5414 23850 5466
rect 23902 5414 23914 5466
rect 23966 5414 23978 5466
rect 24030 5414 26864 5466
rect 1104 5392 26864 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 4571 5324 5365 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 5353 5321 5365 5324
rect 5399 5352 5411 5355
rect 8202 5352 8208 5364
rect 5399 5324 8208 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 8297 5355 8355 5361
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 9030 5352 9036 5364
rect 8343 5324 9036 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 14090 5352 14096 5364
rect 13556 5324 14096 5352
rect 7926 5244 7932 5296
rect 7984 5284 7990 5296
rect 13262 5284 13268 5296
rect 7984 5256 13268 5284
rect 7984 5244 7990 5256
rect 13262 5244 13268 5256
rect 13320 5244 13326 5296
rect 4430 5176 4436 5228
rect 4488 5176 4494 5228
rect 5258 5176 5264 5228
rect 5316 5176 5322 5228
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 6052 5188 7665 5216
rect 6052 5176 6058 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7801 5219 7859 5225
rect 7801 5185 7813 5219
rect 7847 5216 7859 5219
rect 8021 5219 8079 5225
rect 7847 5185 7880 5216
rect 7801 5179 7880 5185
rect 8021 5185 8033 5219
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 4614 5108 4620 5160
rect 4672 5108 4678 5160
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5224 5120 5457 5148
rect 5224 5108 5230 5120
rect 5445 5117 5457 5120
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 7852 5080 7880 5179
rect 8036 5148 8064 5179
rect 8110 5176 8116 5228
rect 8168 5225 8174 5228
rect 8168 5216 8176 5225
rect 8168 5188 8213 5216
rect 8168 5179 8176 5188
rect 8168 5176 8174 5179
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9824 5188 9965 5216
rect 9824 5176 9830 5188
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 13170 5176 13176 5228
rect 13228 5176 13234 5228
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 13556 5216 13584 5324
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 15013 5355 15071 5361
rect 15013 5352 15025 5355
rect 14516 5324 15025 5352
rect 14516 5312 14522 5324
rect 15013 5321 15025 5324
rect 15059 5321 15071 5355
rect 15013 5315 15071 5321
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 16448 5324 16497 5352
rect 16448 5312 16454 5324
rect 16485 5321 16497 5324
rect 16531 5321 16543 5355
rect 16485 5315 16543 5321
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 15372 5287 15430 5293
rect 13648 5256 14872 5284
rect 13648 5228 13676 5256
rect 13403 5188 13584 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 13889 5219 13947 5225
rect 13889 5216 13901 5219
rect 13740 5188 13901 5216
rect 8294 5148 8300 5160
rect 8036 5120 8300 5148
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 10045 5151 10103 5157
rect 10045 5148 10057 5151
rect 9456 5120 10057 5148
rect 9456 5108 9462 5120
rect 10045 5117 10057 5120
rect 10091 5117 10103 5151
rect 10045 5111 10103 5117
rect 10137 5151 10195 5157
rect 10137 5117 10149 5151
rect 10183 5148 10195 5151
rect 13078 5148 13084 5160
rect 10183 5120 13084 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 8202 5080 8208 5092
rect 7852 5052 8208 5080
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 10152 5080 10180 5111
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13740 5148 13768 5188
rect 13889 5185 13901 5188
rect 13935 5185 13947 5219
rect 13889 5179 13947 5185
rect 14844 5160 14872 5256
rect 15372 5253 15384 5287
rect 15418 5284 15430 5287
rect 16684 5284 16712 5315
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 18472 5324 19748 5352
rect 18472 5312 18478 5324
rect 15418 5256 16712 5284
rect 18049 5287 18107 5293
rect 15418 5253 15430 5256
rect 15372 5247 15430 5253
rect 18049 5253 18061 5287
rect 18095 5284 18107 5287
rect 19334 5284 19340 5296
rect 18095 5256 19340 5284
rect 18095 5253 18107 5256
rect 18049 5247 18107 5253
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 19720 5293 19748 5324
rect 19705 5287 19763 5293
rect 19705 5253 19717 5287
rect 19751 5253 19763 5287
rect 21082 5284 21088 5296
rect 19705 5247 19763 5253
rect 20180 5256 21088 5284
rect 16850 5176 16856 5228
rect 16908 5176 16914 5228
rect 17310 5176 17316 5228
rect 17368 5216 17374 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 17368 5188 18245 5216
rect 17368 5176 17374 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18748 5188 18797 5216
rect 18748 5176 18754 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 18966 5176 18972 5228
rect 19024 5176 19030 5228
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5216 19303 5219
rect 20180 5216 20208 5256
rect 21082 5244 21088 5256
rect 21140 5244 21146 5296
rect 19291 5188 20208 5216
rect 20257 5219 20315 5225
rect 19291 5185 19303 5188
rect 19245 5179 19303 5185
rect 20257 5185 20269 5219
rect 20303 5216 20315 5219
rect 20346 5216 20352 5228
rect 20303 5188 20352 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 20346 5176 20352 5188
rect 20404 5176 20410 5228
rect 20438 5176 20444 5228
rect 20496 5176 20502 5228
rect 20714 5176 20720 5228
rect 20772 5176 20778 5228
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 20864 5188 21128 5216
rect 20864 5176 20870 5188
rect 13556 5120 13768 5148
rect 13556 5089 13584 5120
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15105 5151 15163 5157
rect 15105 5148 15117 5151
rect 14884 5120 15117 5148
rect 14884 5108 14890 5120
rect 15105 5117 15117 5120
rect 15151 5117 15163 5151
rect 15105 5111 15163 5117
rect 19153 5151 19211 5157
rect 19153 5117 19165 5151
rect 19199 5117 19211 5151
rect 19153 5111 19211 5117
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5117 19671 5151
rect 19613 5111 19671 5117
rect 8864 5052 10180 5080
rect 13541 5083 13599 5089
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 4028 4984 4077 5012
rect 4028 4972 4034 4984
rect 4065 4981 4077 4984
rect 4111 4981 4123 5015
rect 4065 4975 4123 4981
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4893 5015 4951 5021
rect 4893 5012 4905 5015
rect 4764 4984 4905 5012
rect 4764 4972 4770 4984
rect 4893 4981 4905 4984
rect 4939 4981 4951 5015
rect 4893 4975 4951 4981
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8864 5012 8892 5052
rect 13541 5049 13553 5083
rect 13587 5049 13599 5083
rect 13541 5043 13599 5049
rect 18782 5040 18788 5092
rect 18840 5080 18846 5092
rect 19168 5080 19196 5111
rect 18840 5052 19196 5080
rect 19628 5080 19656 5111
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20456 5148 20484 5176
rect 20036 5120 20484 5148
rect 20901 5151 20959 5157
rect 20036 5108 20042 5120
rect 20901 5117 20913 5151
rect 20947 5148 20959 5151
rect 20990 5148 20996 5160
rect 20947 5120 20996 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 21100 5157 21128 5188
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 20162 5080 20168 5092
rect 19628 5052 20168 5080
rect 18840 5040 18846 5052
rect 7524 4984 8892 5012
rect 7524 4972 7530 4984
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 8996 4984 9597 5012
rect 8996 4972 9002 4984
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 12986 4972 12992 5024
rect 13044 4972 13050 5024
rect 17773 5015 17831 5021
rect 17773 4981 17785 5015
rect 17819 5012 17831 5015
rect 19628 5012 19656 5052
rect 20162 5040 20168 5052
rect 20220 5080 20226 5092
rect 20806 5080 20812 5092
rect 20220 5052 20812 5080
rect 20220 5040 20226 5052
rect 20806 5040 20812 5052
rect 20864 5040 20870 5092
rect 17819 4984 19656 5012
rect 17819 4981 17831 4984
rect 17773 4975 17831 4981
rect 1104 4922 26864 4944
rect 1104 4870 2918 4922
rect 2970 4870 2982 4922
rect 3034 4870 3046 4922
rect 3098 4870 3110 4922
rect 3162 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 6918 4922
rect 6970 4870 6982 4922
rect 7034 4870 7046 4922
rect 7098 4870 7110 4922
rect 7162 4870 7174 4922
rect 7226 4870 7238 4922
rect 7290 4870 10918 4922
rect 10970 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 11238 4922
rect 11290 4870 14918 4922
rect 14970 4870 14982 4922
rect 15034 4870 15046 4922
rect 15098 4870 15110 4922
rect 15162 4870 15174 4922
rect 15226 4870 15238 4922
rect 15290 4870 18918 4922
rect 18970 4870 18982 4922
rect 19034 4870 19046 4922
rect 19098 4870 19110 4922
rect 19162 4870 19174 4922
rect 19226 4870 19238 4922
rect 19290 4870 22918 4922
rect 22970 4870 22982 4922
rect 23034 4870 23046 4922
rect 23098 4870 23110 4922
rect 23162 4870 23174 4922
rect 23226 4870 23238 4922
rect 23290 4870 26864 4922
rect 1104 4848 26864 4870
rect 5994 4768 6000 4820
rect 6052 4768 6058 4820
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 6917 4811 6975 4817
rect 6917 4808 6929 4811
rect 6604 4780 6929 4808
rect 6604 4768 6610 4780
rect 6917 4777 6929 4780
rect 6963 4777 6975 4811
rect 6917 4771 6975 4777
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9272 4780 9413 4808
rect 9272 4768 9278 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 9600 4780 14688 4808
rect 5626 4700 5632 4752
rect 5684 4740 5690 4752
rect 5684 4712 5856 4740
rect 5684 4700 5690 4712
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5316 4644 5764 4672
rect 5316 4632 5322 4644
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 4430 4496 4436 4548
rect 4488 4536 4494 4548
rect 5460 4536 5488 4567
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5736 4613 5764 4644
rect 5828 4613 5856 4712
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 7616 4712 8064 4740
rect 7616 4700 7622 4712
rect 7926 4672 7932 4684
rect 6564 4644 7932 4672
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5592 4576 5641 4604
rect 5592 4564 5598 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 6564 4613 6592 4644
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 8036 4681 8064 4712
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4641 8079 4675
rect 9600 4672 9628 4780
rect 10597 4743 10655 4749
rect 10597 4709 10609 4743
rect 10643 4740 10655 4743
rect 11146 4740 11152 4752
rect 10643 4712 11152 4740
rect 10643 4709 10655 4712
rect 10597 4703 10655 4709
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 13909 4743 13967 4749
rect 13909 4740 13921 4743
rect 13872 4712 13921 4740
rect 13872 4700 13878 4712
rect 13909 4709 13921 4712
rect 13955 4709 13967 4743
rect 14660 4740 14688 4780
rect 14734 4768 14740 4820
rect 14792 4768 14798 4820
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 17218 4808 17224 4820
rect 16715 4780 17224 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 20346 4808 20352 4820
rect 19852 4780 20352 4808
rect 19852 4768 19858 4780
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 20530 4768 20536 4820
rect 20588 4808 20594 4820
rect 22094 4808 22100 4820
rect 20588 4780 22100 4808
rect 20588 4768 20594 4780
rect 22094 4768 22100 4780
rect 22152 4768 22158 4820
rect 14660 4712 14964 4740
rect 13909 4703 13967 4709
rect 14936 4684 14964 4712
rect 18506 4700 18512 4752
rect 18564 4740 18570 4752
rect 18564 4712 20760 4740
rect 18564 4700 18570 4712
rect 8021 4635 8079 4641
rect 9048 4644 9628 4672
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 5960 4576 6377 4604
rect 5960 4564 5966 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 9048 4604 9076 4644
rect 6779 4576 9076 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 9122 4564 9128 4616
rect 9180 4564 9186 4616
rect 9600 4613 9628 4644
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10318 4672 10324 4684
rect 10091 4644 10324 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 10744 4644 11284 4672
rect 10744 4632 10750 4644
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 9766 4564 9772 4616
rect 9824 4564 9830 4616
rect 11256 4613 11284 4644
rect 14918 4632 14924 4684
rect 14976 4672 14982 4684
rect 18322 4672 18328 4684
rect 14976 4644 18328 4672
rect 14976 4632 14982 4644
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 13630 4604 13636 4616
rect 12575 4576 13636 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 4488 4508 5488 4536
rect 4488 4496 4494 4508
rect 6638 4496 6644 4548
rect 6696 4496 6702 4548
rect 7837 4539 7895 4545
rect 7837 4505 7849 4539
rect 7883 4536 7895 4539
rect 8294 4536 8300 4548
rect 7883 4508 8300 4536
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 8294 4496 8300 4508
rect 8352 4496 8358 4548
rect 9398 4536 9404 4548
rect 8404 4508 9404 4536
rect 8404 4480 8432 4508
rect 9398 4496 9404 4508
rect 9456 4536 9462 4548
rect 10137 4539 10195 4545
rect 10137 4536 10149 4539
rect 9456 4508 10149 4536
rect 9456 4496 9462 4508
rect 10137 4505 10149 4508
rect 10183 4505 10195 4539
rect 10778 4536 10784 4548
rect 10137 4499 10195 4505
rect 10244 4508 10784 4536
rect 10244 4480 10272 4508
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 2866 4428 2872 4480
rect 2924 4468 2930 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 2924 4440 3801 4468
rect 2924 4428 2930 4440
rect 3789 4437 3801 4440
rect 3835 4437 3847 4471
rect 3789 4431 3847 4437
rect 4522 4428 4528 4480
rect 4580 4428 4586 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 7156 4440 7481 4468
rect 7156 4428 7162 4440
rect 7469 4437 7481 4440
rect 7515 4437 7527 4471
rect 7469 4431 7527 4437
rect 7929 4471 7987 4477
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8386 4468 8392 4480
rect 7975 4440 8392 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9306 4428 9312 4480
rect 9364 4428 9370 4480
rect 10226 4428 10232 4480
rect 10284 4428 10290 4480
rect 10594 4428 10600 4480
rect 10652 4468 10658 4480
rect 10689 4471 10747 4477
rect 10689 4468 10701 4471
rect 10652 4440 10701 4468
rect 10652 4428 10658 4440
rect 10689 4437 10701 4440
rect 10735 4437 10747 4471
rect 10888 4468 10916 4567
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 14090 4564 14096 4616
rect 14148 4564 14154 4616
rect 14186 4607 14244 4613
rect 14186 4573 14198 4607
rect 14232 4573 14244 4607
rect 14186 4567 14244 4573
rect 10962 4496 10968 4548
rect 11020 4496 11026 4548
rect 11057 4539 11115 4545
rect 11057 4505 11069 4539
rect 11103 4536 11115 4539
rect 12796 4539 12854 4545
rect 11103 4508 12434 4536
rect 11103 4505 11115 4508
rect 11057 4499 11115 4505
rect 11330 4468 11336 4480
rect 10888 4440 11336 4468
rect 10689 4431 10747 4437
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 12406 4468 12434 4508
rect 12796 4505 12808 4539
rect 12842 4536 12854 4539
rect 12986 4536 12992 4548
rect 12842 4508 12992 4536
rect 12842 4505 12854 4508
rect 12796 4499 12854 4505
rect 12986 4496 12992 4508
rect 13044 4496 13050 4548
rect 13906 4496 13912 4548
rect 13964 4536 13970 4548
rect 14200 4536 14228 4567
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 14642 4613 14648 4616
rect 14599 4607 14648 4613
rect 14599 4573 14611 4607
rect 14645 4573 14648 4607
rect 14599 4567 14648 4573
rect 14642 4564 14648 4567
rect 14700 4564 14706 4616
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 17052 4613 17080 4644
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 20732 4681 20760 4712
rect 20717 4675 20775 4681
rect 19444 4644 20576 4672
rect 19444 4616 19472 4644
rect 16807 4607 16865 4613
rect 16807 4604 16819 4607
rect 16632 4576 16819 4604
rect 16632 4564 16638 4576
rect 16807 4573 16819 4576
rect 16853 4573 16865 4607
rect 16807 4567 16865 4573
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4573 17095 4607
rect 17037 4567 17095 4573
rect 17220 4607 17278 4613
rect 17220 4573 17232 4607
rect 17266 4573 17278 4607
rect 17220 4567 17278 4573
rect 13964 4508 14228 4536
rect 14369 4539 14427 4545
rect 13964 4496 13970 4508
rect 14369 4505 14381 4539
rect 14415 4505 14427 4539
rect 14369 4499 14427 4505
rect 14384 4468 14412 4499
rect 16390 4496 16396 4548
rect 16448 4536 16454 4548
rect 16945 4539 17003 4545
rect 16945 4536 16957 4539
rect 16448 4508 16957 4536
rect 16448 4496 16454 4508
rect 16945 4505 16957 4508
rect 16991 4505 17003 4539
rect 17236 4536 17264 4567
rect 17310 4564 17316 4616
rect 17368 4564 17374 4616
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4604 19027 4607
rect 19426 4604 19432 4616
rect 19015 4576 19432 4604
rect 19015 4573 19027 4576
rect 18969 4567 19027 4573
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 19794 4564 19800 4616
rect 19852 4564 19858 4616
rect 19978 4564 19984 4616
rect 20036 4564 20042 4616
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 17402 4536 17408 4548
rect 17236 4508 17408 4536
rect 16945 4499 17003 4505
rect 17402 4496 17408 4508
rect 17460 4496 17466 4548
rect 18782 4496 18788 4548
rect 18840 4536 18846 4548
rect 18877 4539 18935 4545
rect 18877 4536 18889 4539
rect 18840 4508 18889 4536
rect 18840 4496 18846 4508
rect 18877 4505 18889 4508
rect 18923 4536 18935 4539
rect 20180 4536 20208 4567
rect 20254 4564 20260 4616
rect 20312 4564 20318 4616
rect 20548 4548 20576 4644
rect 20717 4641 20729 4675
rect 20763 4672 20775 4675
rect 20763 4644 22416 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 20806 4604 20812 4616
rect 20671 4576 20812 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 20901 4607 20959 4613
rect 20901 4573 20913 4607
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 18923 4508 20208 4536
rect 18923 4505 18935 4508
rect 18877 4499 18935 4505
rect 20530 4496 20536 4548
rect 20588 4536 20594 4548
rect 20916 4536 20944 4567
rect 21910 4564 21916 4616
rect 21968 4564 21974 4616
rect 22186 4564 22192 4616
rect 22244 4564 22250 4616
rect 22388 4613 22416 4644
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 22465 4607 22523 4613
rect 22465 4573 22477 4607
rect 22511 4604 22523 4607
rect 22646 4604 22652 4616
rect 22511 4576 22652 4604
rect 22511 4573 22523 4576
rect 22465 4567 22523 4573
rect 20588 4508 20944 4536
rect 22388 4536 22416 4567
rect 22646 4564 22652 4576
rect 22704 4564 22710 4616
rect 23753 4607 23811 4613
rect 23753 4573 23765 4607
rect 23799 4604 23811 4607
rect 24394 4604 24400 4616
rect 23799 4576 24400 4604
rect 23799 4573 23811 4576
rect 23753 4567 23811 4573
rect 24394 4564 24400 4576
rect 24452 4564 24458 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 25222 4604 25228 4616
rect 24627 4576 25228 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 24210 4536 24216 4548
rect 22388 4508 24216 4536
rect 20588 4496 20594 4508
rect 24210 4496 24216 4508
rect 24268 4496 24274 4548
rect 17862 4468 17868 4480
rect 12406 4440 17868 4468
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 19521 4471 19579 4477
rect 19521 4437 19533 4471
rect 19567 4468 19579 4471
rect 20622 4468 20628 4480
rect 19567 4440 20628 4468
rect 19567 4437 19579 4440
rect 19521 4431 19579 4437
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 21082 4428 21088 4480
rect 21140 4428 21146 4480
rect 21729 4471 21787 4477
rect 21729 4437 21741 4471
rect 21775 4468 21787 4471
rect 22094 4468 22100 4480
rect 21775 4440 22100 4468
rect 21775 4437 21787 4440
rect 21729 4431 21787 4437
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 22554 4428 22560 4480
rect 22612 4428 22618 4480
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 23569 4471 23627 4477
rect 23569 4468 23581 4471
rect 23532 4440 23581 4468
rect 23532 4428 23538 4440
rect 23569 4437 23581 4440
rect 23615 4437 23627 4471
rect 23569 4431 23627 4437
rect 24394 4428 24400 4480
rect 24452 4428 24458 4480
rect 1104 4378 26864 4400
rect 1104 4326 3658 4378
rect 3710 4326 3722 4378
rect 3774 4326 3786 4378
rect 3838 4326 3850 4378
rect 3902 4326 3914 4378
rect 3966 4326 3978 4378
rect 4030 4326 7658 4378
rect 7710 4326 7722 4378
rect 7774 4326 7786 4378
rect 7838 4326 7850 4378
rect 7902 4326 7914 4378
rect 7966 4326 7978 4378
rect 8030 4326 11658 4378
rect 11710 4326 11722 4378
rect 11774 4326 11786 4378
rect 11838 4326 11850 4378
rect 11902 4326 11914 4378
rect 11966 4326 11978 4378
rect 12030 4326 15658 4378
rect 15710 4326 15722 4378
rect 15774 4326 15786 4378
rect 15838 4326 15850 4378
rect 15902 4326 15914 4378
rect 15966 4326 15978 4378
rect 16030 4326 19658 4378
rect 19710 4326 19722 4378
rect 19774 4326 19786 4378
rect 19838 4326 19850 4378
rect 19902 4326 19914 4378
rect 19966 4326 19978 4378
rect 20030 4326 23658 4378
rect 23710 4326 23722 4378
rect 23774 4326 23786 4378
rect 23838 4326 23850 4378
rect 23902 4326 23914 4378
rect 23966 4326 23978 4378
rect 24030 4326 26864 4378
rect 1104 4304 26864 4326
rect 5258 4224 5264 4276
rect 5316 4264 5322 4276
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 5316 4236 5457 4264
rect 5316 4224 5322 4236
rect 5445 4233 5457 4236
rect 5491 4233 5503 4267
rect 5445 4227 5503 4233
rect 6825 4267 6883 4273
rect 6825 4233 6837 4267
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 2866 4205 2872 4208
rect 2860 4159 2872 4205
rect 2924 4196 2930 4208
rect 4332 4199 4390 4205
rect 2924 4168 2960 4196
rect 2866 4156 2872 4159
rect 2924 4156 2930 4168
rect 4332 4165 4344 4199
rect 4378 4196 4390 4199
rect 4522 4196 4528 4208
rect 4378 4168 4528 4196
rect 4378 4165 4390 4168
rect 4332 4159 4390 4165
rect 4522 4156 4528 4168
rect 4580 4156 4586 4208
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2004 4100 2605 4128
rect 2004 4088 2010 4100
rect 2593 4097 2605 4100
rect 2639 4128 2651 4131
rect 4065 4131 4123 4137
rect 4065 4128 4077 4131
rect 2639 4100 4077 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 4065 4097 4077 4100
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6362 4128 6368 4140
rect 5859 4100 6368 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6840 4128 6868 4227
rect 8294 4224 8300 4276
rect 8352 4224 8358 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 9401 4267 9459 4273
rect 9401 4264 9413 4267
rect 9180 4236 9413 4264
rect 9180 4224 9186 4236
rect 9401 4233 9413 4236
rect 9447 4233 9459 4267
rect 10686 4264 10692 4276
rect 9401 4227 9459 4233
rect 10336 4236 10692 4264
rect 9033 4199 9091 4205
rect 9033 4165 9045 4199
rect 9079 4196 9091 4199
rect 10336 4196 10364 4236
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 13081 4267 13139 4273
rect 13081 4233 13093 4267
rect 13127 4264 13139 4267
rect 13170 4264 13176 4276
rect 13127 4236 13176 4264
rect 13127 4233 13139 4236
rect 13081 4227 13139 4233
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 13449 4267 13507 4273
rect 13449 4233 13461 4267
rect 13495 4264 13507 4267
rect 13814 4264 13820 4276
rect 13495 4236 13820 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 13909 4267 13967 4273
rect 13909 4233 13921 4267
rect 13955 4264 13967 4267
rect 14090 4264 14096 4276
rect 13955 4236 14096 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 16114 4224 16120 4276
rect 16172 4224 16178 4276
rect 17310 4224 17316 4276
rect 17368 4264 17374 4276
rect 17497 4267 17555 4273
rect 17497 4264 17509 4267
rect 17368 4236 17509 4264
rect 17368 4224 17374 4236
rect 17497 4233 17509 4236
rect 17543 4233 17555 4267
rect 17497 4227 17555 4233
rect 17862 4224 17868 4276
rect 17920 4264 17926 4276
rect 18138 4264 18144 4276
rect 17920 4236 18144 4264
rect 17920 4224 17926 4236
rect 18138 4224 18144 4236
rect 18196 4224 18202 4276
rect 20070 4224 20076 4276
rect 20128 4224 20134 4276
rect 9079 4168 10364 4196
rect 10428 4168 10916 4196
rect 9079 4165 9091 4168
rect 9033 4159 9091 4165
rect 7173 4131 7231 4137
rect 7173 4128 7185 4131
rect 6687 4100 6776 4128
rect 6840 4100 7185 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 3973 3927 4031 3933
rect 3973 3893 3985 3927
rect 4019 3924 4031 3927
rect 4430 3924 4436 3936
rect 4019 3896 4436 3924
rect 4019 3893 4031 3896
rect 3973 3887 4031 3893
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 5626 3884 5632 3936
rect 5684 3884 5690 3936
rect 6748 3924 6776 4100
rect 7173 4097 7185 4100
rect 7219 4097 7231 4131
rect 7173 4091 7231 4097
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8444 4100 8953 4128
rect 8444 4088 8450 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 10428 4128 10456 4168
rect 9548 4100 10456 4128
rect 9548 4088 9554 4100
rect 10594 4088 10600 4140
rect 10652 4137 10658 4140
rect 10888 4137 10916 4168
rect 13262 4156 13268 4208
rect 13320 4196 13326 4208
rect 14277 4199 14335 4205
rect 14277 4196 14289 4199
rect 13320 4168 14289 4196
rect 13320 4156 13326 4168
rect 14277 4165 14289 4168
rect 14323 4196 14335 4199
rect 16298 4196 16304 4208
rect 14323 4168 16304 4196
rect 14323 4165 14335 4168
rect 14277 4159 14335 4165
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 16960 4168 18000 4196
rect 10652 4128 10664 4137
rect 10873 4131 10931 4137
rect 10652 4100 10697 4128
rect 10652 4091 10664 4100
rect 10873 4097 10885 4131
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 10652 4088 10658 4091
rect 11146 4088 11152 4140
rect 11204 4088 11210 4140
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4128 12679 4131
rect 13354 4128 13360 4140
rect 12667 4100 13360 4128
rect 12667 4097 12679 4100
rect 12621 4091 12679 4097
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13722 4128 13728 4140
rect 13587 4100 13728 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6880 4032 6929 4060
rect 6880 4020 6886 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 8846 4020 8852 4072
rect 8904 4020 8910 4072
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 11388 4032 13645 4060
rect 11388 4020 11394 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 14108 4060 14136 4091
rect 14182 4088 14188 4140
rect 14240 4088 14246 4140
rect 14458 4088 14464 4140
rect 14516 4088 14522 4140
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4128 16083 4131
rect 16390 4128 16396 4140
rect 16071 4100 16396 4128
rect 16071 4097 16083 4100
rect 16025 4091 16083 4097
rect 16390 4088 16396 4100
rect 16448 4128 16454 4140
rect 16960 4128 16988 4168
rect 16448 4100 16988 4128
rect 17037 4131 17095 4137
rect 16448 4088 16454 4100
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17402 4128 17408 4140
rect 17083 4100 17408 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17552 4100 17693 4128
rect 17552 4088 17558 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 14918 4060 14924 4072
rect 14108 4032 14924 4060
rect 13633 4023 13691 4029
rect 13648 3992 13676 4023
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 15028 4032 16313 4060
rect 15028 3992 15056 4032
rect 16301 4029 16313 4032
rect 16347 4060 16359 4063
rect 16666 4060 16672 4072
rect 16347 4032 16672 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17788 4060 17816 4091
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 17972 4128 18000 4168
rect 18690 4156 18696 4208
rect 18748 4196 18754 4208
rect 21082 4196 21088 4208
rect 18748 4168 19104 4196
rect 18748 4156 18754 4168
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17972 4100 18061 4128
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 18598 4088 18604 4140
rect 18656 4128 18662 4140
rect 19076 4137 19104 4168
rect 19720 4168 21088 4196
rect 18969 4131 19027 4137
rect 18969 4128 18981 4131
rect 18656 4100 18981 4128
rect 18656 4088 18662 4100
rect 18969 4097 18981 4100
rect 19015 4097 19027 4131
rect 18969 4091 19027 4097
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 19518 4088 19524 4140
rect 19576 4088 19582 4140
rect 19720 4137 19748 4168
rect 21082 4156 21088 4168
rect 21140 4156 21146 4208
rect 22094 4156 22100 4208
rect 22152 4156 22158 4208
rect 22554 4156 22560 4208
rect 22612 4156 22618 4208
rect 24210 4196 24216 4208
rect 23860 4168 24216 4196
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 19978 4128 19984 4140
rect 19935 4100 19984 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 18322 4060 18328 4072
rect 17788 4032 18328 4060
rect 17313 4023 17371 4029
rect 13648 3964 15056 3992
rect 16206 3952 16212 4004
rect 16264 3992 16270 4004
rect 17144 3992 17172 4023
rect 16264 3964 17172 3992
rect 17328 3992 17356 4023
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 17328 3964 18000 3992
rect 16264 3952 16270 3964
rect 17972 3936 18000 3964
rect 18506 3952 18512 4004
rect 18564 3992 18570 4004
rect 20088 3992 20116 4091
rect 20530 4088 20536 4140
rect 20588 4088 20594 4140
rect 23860 4137 23888 4168
rect 24210 4156 24216 4168
rect 24268 4156 24274 4208
rect 24305 4199 24363 4205
rect 24305 4165 24317 4199
rect 24351 4196 24363 4199
rect 24394 4196 24400 4208
rect 24351 4168 24400 4196
rect 24351 4165 24363 4168
rect 24305 4159 24363 4165
rect 24394 4156 24400 4168
rect 24452 4156 24458 4208
rect 24946 4156 24952 4208
rect 25004 4156 25010 4208
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 26053 4131 26111 4137
rect 26053 4128 26065 4131
rect 25740 4100 26065 4128
rect 25740 4088 25746 4100
rect 26053 4097 26065 4100
rect 26099 4097 26111 4131
rect 26053 4091 26111 4097
rect 21821 4063 21879 4069
rect 21821 4029 21833 4063
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 24029 4063 24087 4069
rect 24029 4029 24041 4063
rect 24075 4029 24087 4063
rect 24029 4023 24087 4029
rect 18564 3964 20116 3992
rect 18564 3952 18570 3964
rect 7098 3924 7104 3936
rect 6748 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 9493 3927 9551 3933
rect 9493 3893 9505 3927
rect 9539 3924 9551 3927
rect 10226 3924 10232 3936
rect 9539 3896 10232 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 10965 3927 11023 3933
rect 10965 3924 10977 3927
rect 10652 3896 10977 3924
rect 10652 3884 10658 3896
rect 10965 3893 10977 3896
rect 11011 3893 11023 3927
rect 10965 3887 11023 3893
rect 12434 3884 12440 3936
rect 12492 3884 12498 3936
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15620 3896 15669 3924
rect 15620 3884 15626 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 16172 3896 16681 3924
rect 16172 3884 16178 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18601 3927 18659 3933
rect 18601 3924 18613 3927
rect 18012 3896 18613 3924
rect 18012 3884 18018 3896
rect 18601 3893 18613 3896
rect 18647 3893 18659 3927
rect 18601 3887 18659 3893
rect 21450 3884 21456 3936
rect 21508 3924 21514 3936
rect 21836 3924 21864 4023
rect 22462 3924 22468 3936
rect 21508 3896 22468 3924
rect 21508 3884 21514 3896
rect 22462 3884 22468 3896
rect 22520 3924 22526 3936
rect 24044 3924 24072 4023
rect 22520 3896 24072 3924
rect 22520 3884 22526 3896
rect 1104 3834 26864 3856
rect 1104 3782 2918 3834
rect 2970 3782 2982 3834
rect 3034 3782 3046 3834
rect 3098 3782 3110 3834
rect 3162 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 6918 3834
rect 6970 3782 6982 3834
rect 7034 3782 7046 3834
rect 7098 3782 7110 3834
rect 7162 3782 7174 3834
rect 7226 3782 7238 3834
rect 7290 3782 10918 3834
rect 10970 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 11238 3834
rect 11290 3782 14918 3834
rect 14970 3782 14982 3834
rect 15034 3782 15046 3834
rect 15098 3782 15110 3834
rect 15162 3782 15174 3834
rect 15226 3782 15238 3834
rect 15290 3782 18918 3834
rect 18970 3782 18982 3834
rect 19034 3782 19046 3834
rect 19098 3782 19110 3834
rect 19162 3782 19174 3834
rect 19226 3782 19238 3834
rect 19290 3782 22918 3834
rect 22970 3782 22982 3834
rect 23034 3782 23046 3834
rect 23098 3782 23110 3834
rect 23162 3782 23174 3834
rect 23226 3782 23238 3834
rect 23290 3782 26864 3834
rect 1104 3760 26864 3782
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 6638 3720 6644 3732
rect 6595 3692 6644 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 8202 3680 8208 3732
rect 8260 3680 8266 3732
rect 9490 3720 9496 3732
rect 9232 3692 9496 3720
rect 9232 3596 9260 3692
rect 9490 3680 9496 3692
rect 9548 3720 9554 3732
rect 13541 3723 13599 3729
rect 9548 3692 12204 3720
rect 9548 3680 9554 3692
rect 10597 3655 10655 3661
rect 10597 3621 10609 3655
rect 10643 3652 10655 3655
rect 10686 3652 10692 3664
rect 10643 3624 10692 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 9214 3544 9220 3596
rect 9272 3544 9278 3596
rect 12066 3544 12072 3596
rect 12124 3584 12130 3596
rect 12176 3593 12204 3692
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 14182 3720 14188 3732
rect 13587 3692 14188 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 15028 3692 15976 3720
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 12124 3556 12173 3584
rect 12124 3544 12130 3556
rect 12161 3553 12173 3556
rect 12207 3553 12219 3587
rect 12161 3547 12219 3553
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 13780 3556 14565 3584
rect 13780 3544 13786 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 15028 3584 15056 3692
rect 15948 3652 15976 3692
rect 16390 3680 16396 3732
rect 16448 3680 16454 3732
rect 16758 3720 16764 3732
rect 16500 3692 16764 3720
rect 16500 3652 16528 3692
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17460 3692 17877 3720
rect 17460 3680 17466 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 21910 3720 21916 3732
rect 17865 3683 17923 3689
rect 21284 3692 21916 3720
rect 15948 3624 16528 3652
rect 18693 3655 18751 3661
rect 18693 3621 18705 3655
rect 18739 3621 18751 3655
rect 18693 3615 18751 3621
rect 14792 3556 15056 3584
rect 18141 3587 18199 3593
rect 14792 3544 14798 3556
rect 18141 3553 18153 3587
rect 18187 3584 18199 3587
rect 18414 3584 18420 3596
rect 18187 3556 18420 3584
rect 18187 3553 18199 3556
rect 18141 3547 18199 3553
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 4706 3476 4712 3528
rect 4764 3476 4770 3528
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 6822 3516 6828 3528
rect 5224 3488 6828 3516
rect 5224 3476 5230 3488
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 8938 3476 8944 3528
rect 8996 3476 9002 3528
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 12434 3525 12440 3528
rect 9473 3519 9531 3525
rect 9473 3516 9485 3519
rect 9364 3488 9485 3516
rect 9364 3476 9370 3488
rect 9473 3485 9485 3488
rect 9519 3485 9531 3519
rect 9473 3479 9531 3485
rect 11885 3519 11943 3525
rect 11885 3485 11897 3519
rect 11931 3485 11943 3519
rect 11885 3479 11943 3485
rect 12428 3479 12440 3525
rect 12492 3516 12498 3528
rect 12492 3488 12528 3516
rect 5436 3451 5494 3457
rect 5436 3417 5448 3451
rect 5482 3448 5494 3451
rect 5626 3448 5632 3460
rect 5482 3420 5632 3448
rect 5482 3417 5494 3420
rect 5436 3411 5494 3417
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 7092 3451 7150 3457
rect 7092 3417 7104 3451
rect 7138 3448 7150 3451
rect 7190 3448 7196 3460
rect 7138 3420 7196 3448
rect 7138 3417 7150 3420
rect 7092 3411 7150 3417
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 8846 3408 8852 3460
rect 8904 3448 8910 3460
rect 11330 3448 11336 3460
rect 8904 3420 11336 3448
rect 8904 3408 8910 3420
rect 11330 3408 11336 3420
rect 11388 3408 11394 3460
rect 11900 3448 11928 3479
rect 12434 3476 12440 3479
rect 12492 3476 12498 3488
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 14458 3516 14464 3528
rect 13320 3488 14464 3516
rect 13320 3476 13326 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14884 3488 15025 3516
rect 14884 3476 14890 3488
rect 15013 3485 15025 3488
rect 15059 3516 15071 3519
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 15059 3488 16497 3516
rect 15059 3485 15071 3488
rect 15013 3479 15071 3485
rect 16485 3485 16497 3488
rect 16531 3485 16543 3519
rect 18708 3516 18736 3615
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3584 21143 3587
rect 21284 3584 21312 3692
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 24946 3680 24952 3732
rect 25004 3680 25010 3732
rect 21131 3556 21312 3584
rect 21361 3587 21419 3593
rect 21131 3553 21143 3556
rect 21085 3547 21143 3553
rect 21361 3553 21373 3587
rect 21407 3584 21419 3587
rect 21729 3587 21787 3593
rect 21729 3584 21741 3587
rect 21407 3556 21741 3584
rect 21407 3553 21419 3556
rect 21361 3547 21419 3553
rect 21729 3553 21741 3556
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 23477 3587 23535 3593
rect 23477 3584 23489 3587
rect 22796 3556 23489 3584
rect 22796 3544 22802 3556
rect 23477 3553 23489 3556
rect 23523 3553 23535 3587
rect 23477 3547 23535 3553
rect 18969 3519 19027 3525
rect 18969 3516 18981 3519
rect 18708 3488 18981 3516
rect 16485 3479 16543 3485
rect 18969 3485 18981 3488
rect 19015 3485 19027 3519
rect 18969 3479 19027 3485
rect 20993 3519 21051 3525
rect 20993 3485 21005 3519
rect 21039 3485 21051 3519
rect 20993 3479 21051 3485
rect 15280 3451 15338 3457
rect 11900 3420 14136 3448
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 9122 3340 9128 3392
rect 9180 3340 9186 3392
rect 12069 3383 12127 3389
rect 12069 3349 12081 3383
rect 12115 3380 12127 3383
rect 12250 3380 12256 3392
rect 12115 3352 12256 3380
rect 12115 3349 12127 3352
rect 12069 3343 12127 3349
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 14108 3389 14136 3420
rect 15280 3417 15292 3451
rect 15326 3448 15338 3451
rect 15378 3448 15384 3460
rect 15326 3420 15384 3448
rect 15326 3417 15338 3420
rect 15280 3411 15338 3417
rect 15378 3408 15384 3420
rect 15436 3408 15442 3460
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 16730 3451 16788 3457
rect 16730 3448 16742 3451
rect 16356 3420 16742 3448
rect 16356 3408 16362 3420
rect 16730 3417 16742 3420
rect 16776 3417 16788 3451
rect 16730 3411 16788 3417
rect 14093 3383 14151 3389
rect 14093 3349 14105 3383
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 16264 3352 18245 3380
rect 16264 3340 16270 3352
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 18322 3340 18328 3392
rect 18380 3340 18386 3392
rect 18782 3340 18788 3392
rect 18840 3340 18846 3392
rect 21008 3380 21036 3479
rect 21450 3476 21456 3528
rect 21508 3476 21514 3528
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 23072 3488 24593 3516
rect 23072 3476 23078 3488
rect 24581 3485 24593 3488
rect 24627 3516 24639 3519
rect 24857 3519 24915 3525
rect 24857 3516 24869 3519
rect 24627 3488 24869 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 24857 3485 24869 3488
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 22462 3408 22468 3460
rect 22520 3408 22526 3460
rect 22738 3380 22744 3392
rect 21008 3352 22744 3380
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 24486 3340 24492 3392
rect 24544 3340 24550 3392
rect 1104 3290 26864 3312
rect 1104 3238 3658 3290
rect 3710 3238 3722 3290
rect 3774 3238 3786 3290
rect 3838 3238 3850 3290
rect 3902 3238 3914 3290
rect 3966 3238 3978 3290
rect 4030 3238 7658 3290
rect 7710 3238 7722 3290
rect 7774 3238 7786 3290
rect 7838 3238 7850 3290
rect 7902 3238 7914 3290
rect 7966 3238 7978 3290
rect 8030 3238 11658 3290
rect 11710 3238 11722 3290
rect 11774 3238 11786 3290
rect 11838 3238 11850 3290
rect 11902 3238 11914 3290
rect 11966 3238 11978 3290
rect 12030 3238 15658 3290
rect 15710 3238 15722 3290
rect 15774 3238 15786 3290
rect 15838 3238 15850 3290
rect 15902 3238 15914 3290
rect 15966 3238 15978 3290
rect 16030 3238 19658 3290
rect 19710 3238 19722 3290
rect 19774 3238 19786 3290
rect 19838 3238 19850 3290
rect 19902 3238 19914 3290
rect 19966 3238 19978 3290
rect 20030 3238 23658 3290
rect 23710 3238 23722 3290
rect 23774 3238 23786 3290
rect 23838 3238 23850 3290
rect 23902 3238 23914 3290
rect 23966 3238 23978 3290
rect 24030 3238 26864 3290
rect 1104 3216 26864 3238
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 4764 3148 5457 3176
rect 4764 3136 4770 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 5902 3176 5908 3188
rect 5859 3148 5908 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6362 3136 6368 3188
rect 6420 3136 6426 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 6733 3179 6791 3185
rect 6733 3176 6745 3179
rect 6696 3148 6745 3176
rect 6696 3136 6702 3148
rect 6733 3145 6745 3148
rect 6779 3145 6791 3179
rect 6733 3139 6791 3145
rect 7190 3136 7196 3188
rect 7248 3136 7254 3188
rect 7469 3179 7527 3185
rect 7469 3145 7481 3179
rect 7515 3145 7527 3179
rect 7469 3139 7527 3145
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8202 3176 8208 3188
rect 7883 3148 8208 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 5166 3108 5172 3120
rect 3988 3080 5172 3108
rect 3988 3049 4016 3080
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4240 3043 4298 3049
rect 4240 3009 4252 3043
rect 4286 3040 4298 3043
rect 4522 3040 4528 3052
rect 4286 3012 4528 3040
rect 4286 3009 4298 3012
rect 4240 3003 4298 3009
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 6270 3040 6276 3052
rect 5951 3012 6276 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6270 3000 6276 3012
rect 6328 3040 6334 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6328 3012 6837 3040
rect 6328 3000 6334 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7484 3040 7512 3139
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9824 3148 10609 3176
rect 9824 3136 9830 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 13262 3136 13268 3188
rect 13320 3136 13326 3188
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 14182 3176 14188 3188
rect 13771 3148 14188 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 15378 3136 15384 3188
rect 15436 3136 15442 3188
rect 16298 3136 16304 3188
rect 16356 3136 16362 3188
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 18322 3176 18328 3188
rect 17083 3148 18328 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 22462 3136 22468 3188
rect 22520 3176 22526 3188
rect 22557 3179 22615 3185
rect 22557 3176 22569 3179
rect 22520 3148 22569 3176
rect 22520 3136 22526 3148
rect 22557 3145 22569 3148
rect 22603 3145 22615 3179
rect 22557 3139 22615 3145
rect 24302 3136 24308 3188
rect 24360 3176 24366 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 24360 3148 24869 3176
rect 24360 3136 24366 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 9122 3068 9128 3120
rect 9180 3108 9186 3120
rect 9462 3111 9520 3117
rect 9462 3108 9474 3111
rect 9180 3080 9474 3108
rect 9180 3068 9186 3080
rect 9462 3077 9474 3080
rect 9508 3077 9520 3111
rect 12066 3108 12072 3120
rect 9462 3071 9520 3077
rect 11900 3080 12072 3108
rect 7423 3012 7512 3040
rect 7929 3043 7987 3049
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8386 3040 8392 3052
rect 7975 3012 8392 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 9214 3000 9220 3052
rect 9272 3000 9278 3052
rect 11900 3049 11928 3080
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 12250 3068 12256 3120
rect 12308 3068 12314 3120
rect 13078 3068 13084 3120
rect 13136 3108 13142 3120
rect 17954 3108 17960 3120
rect 13136 3080 17960 3108
rect 13136 3068 13142 3080
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 12152 3043 12210 3049
rect 12152 3009 12164 3043
rect 12198 3040 12210 3043
rect 12268 3040 12296 3068
rect 12198 3012 12296 3040
rect 12198 3009 12210 3012
rect 12152 3003 12210 3009
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13780 3012 13829 3040
rect 13780 3000 13786 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 6089 2975 6147 2981
rect 6089 2941 6101 2975
rect 6135 2941 6147 2975
rect 6089 2935 6147 2941
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7466 2972 7472 2984
rect 7055 2944 7472 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 6104 2904 6132 2935
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 14016 2981 14044 3080
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 18172 3111 18230 3117
rect 18172 3077 18184 3111
rect 18218 3108 18230 3111
rect 18782 3108 18788 3120
rect 18218 3080 18788 3108
rect 18218 3077 18230 3080
rect 18172 3071 18230 3077
rect 18782 3068 18788 3080
rect 18840 3068 18846 3120
rect 23385 3111 23443 3117
rect 23385 3077 23397 3111
rect 23431 3108 23443 3111
rect 23474 3108 23480 3120
rect 23431 3080 23480 3108
rect 23431 3077 23443 3080
rect 23385 3071 23443 3077
rect 23474 3068 23480 3080
rect 23532 3068 23538 3120
rect 15562 3000 15568 3052
rect 15620 3000 15626 3052
rect 16114 3000 16120 3052
rect 16172 3000 16178 3052
rect 22465 3043 22523 3049
rect 22465 3009 22477 3043
rect 22511 3040 22523 3043
rect 22646 3040 22652 3052
rect 22511 3012 22652 3040
rect 22511 3009 22523 3012
rect 22465 3003 22523 3009
rect 22646 3000 22652 3012
rect 22704 3040 22710 3052
rect 23014 3040 23020 3052
rect 22704 3012 23020 3040
rect 22704 3000 22710 3012
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 24486 3000 24492 3052
rect 24544 3000 24550 3052
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2941 8171 2975
rect 8113 2935 8171 2941
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2972 18475 2975
rect 21450 2972 21456 2984
rect 18463 2944 21456 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 8128 2904 8156 2935
rect 21450 2932 21456 2944
rect 21508 2972 21514 2984
rect 23109 2975 23167 2981
rect 23109 2972 23121 2975
rect 21508 2944 23121 2972
rect 21508 2932 21514 2944
rect 23109 2941 23121 2944
rect 23155 2941 23167 2975
rect 23109 2935 23167 2941
rect 4908 2876 8156 2904
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 4908 2836 4936 2876
rect 4212 2808 4936 2836
rect 5353 2839 5411 2845
rect 4212 2796 4218 2808
rect 5353 2805 5365 2839
rect 5399 2836 5411 2839
rect 5902 2836 5908 2848
rect 5399 2808 5908 2836
rect 5399 2805 5411 2808
rect 5353 2799 5411 2805
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 8128 2836 8156 2876
rect 14734 2836 14740 2848
rect 8128 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 1104 2746 26864 2768
rect 1104 2694 2918 2746
rect 2970 2694 2982 2746
rect 3034 2694 3046 2746
rect 3098 2694 3110 2746
rect 3162 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 6918 2746
rect 6970 2694 6982 2746
rect 7034 2694 7046 2746
rect 7098 2694 7110 2746
rect 7162 2694 7174 2746
rect 7226 2694 7238 2746
rect 7290 2694 10918 2746
rect 10970 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 11238 2746
rect 11290 2694 14918 2746
rect 14970 2694 14982 2746
rect 15034 2694 15046 2746
rect 15098 2694 15110 2746
rect 15162 2694 15174 2746
rect 15226 2694 15238 2746
rect 15290 2694 18918 2746
rect 18970 2694 18982 2746
rect 19034 2694 19046 2746
rect 19098 2694 19110 2746
rect 19162 2694 19174 2746
rect 19226 2694 19238 2746
rect 19290 2694 22918 2746
rect 22970 2694 22982 2746
rect 23034 2694 23046 2746
rect 23098 2694 23110 2746
rect 23162 2694 23174 2746
rect 23226 2694 23238 2746
rect 23290 2694 26864 2746
rect 1104 2672 26864 2694
rect 5997 2635 6055 2641
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 6270 2632 6276 2644
rect 6043 2604 6276 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 8386 2524 8392 2576
rect 8444 2564 8450 2576
rect 8444 2536 9260 2564
rect 8444 2524 8450 2536
rect 9232 2505 9260 2536
rect 16206 2524 16212 2576
rect 16264 2524 16270 2576
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2465 9275 2499
rect 9217 2459 9275 2465
rect 13265 2499 13323 2505
rect 13265 2465 13277 2499
rect 13311 2496 13323 2499
rect 13630 2496 13636 2508
rect 13311 2468 13636 2496
rect 13311 2465 13323 2468
rect 13265 2459 13323 2465
rect 13630 2456 13636 2468
rect 13688 2456 13694 2508
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 5868 2400 6929 2428
rect 5868 2388 5874 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2428 8263 2431
rect 8386 2428 8392 2440
rect 8251 2400 8392 2428
rect 8251 2397 8263 2400
rect 8205 2391 8263 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8803 2400 8953 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12802 2428 12808 2440
rect 12391 2400 12808 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2428 12955 2431
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12943 2400 13001 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 17221 2431 17279 2437
rect 17221 2428 17233 2431
rect 16172 2400 17233 2428
rect 16172 2388 16178 2400
rect 17221 2397 17233 2400
rect 17267 2397 17279 2431
rect 17221 2391 17279 2397
rect 6089 2363 6147 2369
rect 6089 2329 6101 2363
rect 6135 2360 6147 2363
rect 6365 2363 6423 2369
rect 6365 2360 6377 2363
rect 6135 2332 6377 2360
rect 6135 2329 6147 2332
rect 6089 2323 6147 2329
rect 6365 2329 6377 2332
rect 6411 2329 6423 2363
rect 6365 2323 6423 2329
rect 16393 2363 16451 2369
rect 16393 2329 16405 2363
rect 16439 2360 16451 2363
rect 16669 2363 16727 2369
rect 16669 2360 16681 2363
rect 16439 2332 16681 2360
rect 16439 2329 16451 2332
rect 16393 2323 16451 2329
rect 16669 2329 16681 2332
rect 16715 2329 16727 2363
rect 16669 2323 16727 2329
rect 1104 2202 26864 2224
rect 1104 2150 3658 2202
rect 3710 2150 3722 2202
rect 3774 2150 3786 2202
rect 3838 2150 3850 2202
rect 3902 2150 3914 2202
rect 3966 2150 3978 2202
rect 4030 2150 7658 2202
rect 7710 2150 7722 2202
rect 7774 2150 7786 2202
rect 7838 2150 7850 2202
rect 7902 2150 7914 2202
rect 7966 2150 7978 2202
rect 8030 2150 11658 2202
rect 11710 2150 11722 2202
rect 11774 2150 11786 2202
rect 11838 2150 11850 2202
rect 11902 2150 11914 2202
rect 11966 2150 11978 2202
rect 12030 2150 15658 2202
rect 15710 2150 15722 2202
rect 15774 2150 15786 2202
rect 15838 2150 15850 2202
rect 15902 2150 15914 2202
rect 15966 2150 15978 2202
rect 16030 2150 19658 2202
rect 19710 2150 19722 2202
rect 19774 2150 19786 2202
rect 19838 2150 19850 2202
rect 19902 2150 19914 2202
rect 19966 2150 19978 2202
rect 20030 2150 23658 2202
rect 23710 2150 23722 2202
rect 23774 2150 23786 2202
rect 23838 2150 23850 2202
rect 23902 2150 23914 2202
rect 23966 2150 23978 2202
rect 24030 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 2918 27718 2970 27770
rect 2982 27718 3034 27770
rect 3046 27718 3098 27770
rect 3110 27718 3162 27770
rect 3174 27718 3226 27770
rect 3238 27718 3290 27770
rect 6918 27718 6970 27770
rect 6982 27718 7034 27770
rect 7046 27718 7098 27770
rect 7110 27718 7162 27770
rect 7174 27718 7226 27770
rect 7238 27718 7290 27770
rect 10918 27718 10970 27770
rect 10982 27718 11034 27770
rect 11046 27718 11098 27770
rect 11110 27718 11162 27770
rect 11174 27718 11226 27770
rect 11238 27718 11290 27770
rect 14918 27718 14970 27770
rect 14982 27718 15034 27770
rect 15046 27718 15098 27770
rect 15110 27718 15162 27770
rect 15174 27718 15226 27770
rect 15238 27718 15290 27770
rect 18918 27718 18970 27770
rect 18982 27718 19034 27770
rect 19046 27718 19098 27770
rect 19110 27718 19162 27770
rect 19174 27718 19226 27770
rect 19238 27718 19290 27770
rect 22918 27718 22970 27770
rect 22982 27718 23034 27770
rect 23046 27718 23098 27770
rect 23110 27718 23162 27770
rect 23174 27718 23226 27770
rect 23238 27718 23290 27770
rect 9772 27591 9824 27600
rect 9772 27557 9781 27591
rect 9781 27557 9815 27591
rect 9815 27557 9824 27591
rect 9772 27548 9824 27557
rect 10324 27548 10376 27600
rect 10784 27548 10836 27600
rect 11704 27591 11756 27600
rect 11704 27557 11713 27591
rect 11713 27557 11747 27591
rect 11747 27557 11756 27591
rect 11704 27548 11756 27557
rect 12348 27591 12400 27600
rect 12348 27557 12357 27591
rect 12357 27557 12391 27591
rect 12391 27557 12400 27591
rect 12348 27548 12400 27557
rect 14280 27591 14332 27600
rect 14280 27557 14289 27591
rect 14289 27557 14323 27591
rect 14323 27557 14332 27591
rect 14280 27548 14332 27557
rect 17408 27548 17460 27600
rect 20076 27591 20128 27600
rect 20076 27557 20085 27591
rect 20085 27557 20119 27591
rect 20119 27557 20128 27591
rect 20076 27548 20128 27557
rect 20628 27480 20680 27532
rect 9772 27412 9824 27464
rect 10600 27455 10652 27464
rect 10600 27421 10609 27455
rect 10609 27421 10643 27455
rect 10643 27421 10652 27455
rect 10600 27412 10652 27421
rect 11520 27412 11572 27464
rect 11428 27344 11480 27396
rect 12164 27412 12216 27464
rect 14464 27455 14516 27464
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 17684 27455 17736 27464
rect 17684 27421 17693 27455
rect 17693 27421 17727 27455
rect 17727 27421 17736 27455
rect 17684 27412 17736 27421
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 19524 27412 19576 27464
rect 20076 27412 20128 27464
rect 20536 27412 20588 27464
rect 18696 27276 18748 27328
rect 21088 27276 21140 27328
rect 3658 27174 3710 27226
rect 3722 27174 3774 27226
rect 3786 27174 3838 27226
rect 3850 27174 3902 27226
rect 3914 27174 3966 27226
rect 3978 27174 4030 27226
rect 7658 27174 7710 27226
rect 7722 27174 7774 27226
rect 7786 27174 7838 27226
rect 7850 27174 7902 27226
rect 7914 27174 7966 27226
rect 7978 27174 8030 27226
rect 11658 27174 11710 27226
rect 11722 27174 11774 27226
rect 11786 27174 11838 27226
rect 11850 27174 11902 27226
rect 11914 27174 11966 27226
rect 11978 27174 12030 27226
rect 15658 27174 15710 27226
rect 15722 27174 15774 27226
rect 15786 27174 15838 27226
rect 15850 27174 15902 27226
rect 15914 27174 15966 27226
rect 15978 27174 16030 27226
rect 19658 27174 19710 27226
rect 19722 27174 19774 27226
rect 19786 27174 19838 27226
rect 19850 27174 19902 27226
rect 19914 27174 19966 27226
rect 19978 27174 20030 27226
rect 23658 27174 23710 27226
rect 23722 27174 23774 27226
rect 23786 27174 23838 27226
rect 23850 27174 23902 27226
rect 23914 27174 23966 27226
rect 23978 27174 24030 27226
rect 4988 26979 5040 26988
rect 4988 26945 4997 26979
rect 4997 26945 5031 26979
rect 5031 26945 5040 26979
rect 4988 26936 5040 26945
rect 9772 27072 9824 27124
rect 8760 26936 8812 26988
rect 8392 26911 8444 26920
rect 8392 26877 8401 26911
rect 8401 26877 8435 26911
rect 8435 26877 8444 26911
rect 8392 26868 8444 26877
rect 8576 26911 8628 26920
rect 8576 26877 8585 26911
rect 8585 26877 8619 26911
rect 8619 26877 8628 26911
rect 8576 26868 8628 26877
rect 9312 26868 9364 26920
rect 9680 26800 9732 26852
rect 10232 26979 10284 26988
rect 10232 26945 10241 26979
rect 10241 26945 10275 26979
rect 10275 26945 10284 26979
rect 10232 26936 10284 26945
rect 10784 27004 10836 27056
rect 11060 27072 11112 27124
rect 12532 27004 12584 27056
rect 10692 26979 10744 26988
rect 10692 26945 10701 26979
rect 10701 26945 10735 26979
rect 10735 26945 10744 26979
rect 10692 26936 10744 26945
rect 10876 26979 10928 26988
rect 10876 26945 10885 26979
rect 10885 26945 10919 26979
rect 10919 26945 10928 26979
rect 10876 26936 10928 26945
rect 10600 26868 10652 26920
rect 11888 26868 11940 26920
rect 12992 26979 13044 26988
rect 12992 26945 13001 26979
rect 13001 26945 13035 26979
rect 13035 26945 13044 26979
rect 12992 26936 13044 26945
rect 13544 26979 13596 26988
rect 13544 26945 13553 26979
rect 13553 26945 13587 26979
rect 13587 26945 13596 26979
rect 13544 26936 13596 26945
rect 4804 26775 4856 26784
rect 4804 26741 4813 26775
rect 4813 26741 4847 26775
rect 4847 26741 4856 26775
rect 4804 26732 4856 26741
rect 7656 26775 7708 26784
rect 7656 26741 7665 26775
rect 7665 26741 7699 26775
rect 7699 26741 7708 26775
rect 7656 26732 7708 26741
rect 9220 26732 9272 26784
rect 10508 26732 10560 26784
rect 10784 26800 10836 26852
rect 14832 26936 14884 26988
rect 19432 27072 19484 27124
rect 20904 27072 20956 27124
rect 19524 27004 19576 27056
rect 20352 27004 20404 27056
rect 13820 26868 13872 26920
rect 17224 26979 17276 26988
rect 17224 26945 17233 26979
rect 17233 26945 17267 26979
rect 17267 26945 17276 26979
rect 17224 26936 17276 26945
rect 17592 26936 17644 26988
rect 18604 26936 18656 26988
rect 20812 26936 20864 26988
rect 16580 26868 16632 26920
rect 17408 26868 17460 26920
rect 14464 26800 14516 26852
rect 10968 26732 11020 26784
rect 11336 26732 11388 26784
rect 12716 26732 12768 26784
rect 13360 26775 13412 26784
rect 13360 26741 13369 26775
rect 13369 26741 13403 26775
rect 13403 26741 13412 26775
rect 13360 26732 13412 26741
rect 13912 26732 13964 26784
rect 14648 26775 14700 26784
rect 14648 26741 14657 26775
rect 14657 26741 14691 26775
rect 14691 26741 14700 26775
rect 14648 26732 14700 26741
rect 14740 26732 14792 26784
rect 16488 26732 16540 26784
rect 17500 26800 17552 26852
rect 18788 26911 18840 26920
rect 18788 26877 18797 26911
rect 18797 26877 18831 26911
rect 18831 26877 18840 26911
rect 18788 26868 18840 26877
rect 17224 26732 17276 26784
rect 17408 26775 17460 26784
rect 17408 26741 17417 26775
rect 17417 26741 17451 26775
rect 17451 26741 17460 26775
rect 17408 26732 17460 26741
rect 17868 26732 17920 26784
rect 20076 26732 20128 26784
rect 20260 26732 20312 26784
rect 2918 26630 2970 26682
rect 2982 26630 3034 26682
rect 3046 26630 3098 26682
rect 3110 26630 3162 26682
rect 3174 26630 3226 26682
rect 3238 26630 3290 26682
rect 6918 26630 6970 26682
rect 6982 26630 7034 26682
rect 7046 26630 7098 26682
rect 7110 26630 7162 26682
rect 7174 26630 7226 26682
rect 7238 26630 7290 26682
rect 10918 26630 10970 26682
rect 10982 26630 11034 26682
rect 11046 26630 11098 26682
rect 11110 26630 11162 26682
rect 11174 26630 11226 26682
rect 11238 26630 11290 26682
rect 14918 26630 14970 26682
rect 14982 26630 15034 26682
rect 15046 26630 15098 26682
rect 15110 26630 15162 26682
rect 15174 26630 15226 26682
rect 15238 26630 15290 26682
rect 18918 26630 18970 26682
rect 18982 26630 19034 26682
rect 19046 26630 19098 26682
rect 19110 26630 19162 26682
rect 19174 26630 19226 26682
rect 19238 26630 19290 26682
rect 22918 26630 22970 26682
rect 22982 26630 23034 26682
rect 23046 26630 23098 26682
rect 23110 26630 23162 26682
rect 23174 26630 23226 26682
rect 23238 26630 23290 26682
rect 5080 26528 5132 26580
rect 8760 26571 8812 26580
rect 8760 26537 8769 26571
rect 8769 26537 8803 26571
rect 8803 26537 8812 26571
rect 8760 26528 8812 26537
rect 9036 26528 9088 26580
rect 11888 26571 11940 26580
rect 11888 26537 11897 26571
rect 11897 26537 11931 26571
rect 11931 26537 11940 26571
rect 11888 26528 11940 26537
rect 16672 26528 16724 26580
rect 5448 26392 5500 26444
rect 7012 26392 7064 26444
rect 7196 26392 7248 26444
rect 4068 26367 4120 26376
rect 4068 26333 4077 26367
rect 4077 26333 4111 26367
rect 4111 26333 4120 26367
rect 4068 26324 4120 26333
rect 4436 26367 4488 26376
rect 4436 26333 4445 26367
rect 4445 26333 4479 26367
rect 4479 26333 4488 26367
rect 17592 26503 17644 26512
rect 17592 26469 17601 26503
rect 17601 26469 17635 26503
rect 17635 26469 17644 26503
rect 17592 26460 17644 26469
rect 7380 26435 7432 26444
rect 7380 26401 7389 26435
rect 7389 26401 7423 26435
rect 7423 26401 7432 26435
rect 7380 26392 7432 26401
rect 8576 26392 8628 26444
rect 10416 26392 10468 26444
rect 4436 26324 4488 26333
rect 7656 26367 7708 26376
rect 7656 26333 7690 26367
rect 7690 26333 7708 26367
rect 7656 26324 7708 26333
rect 12256 26324 12308 26376
rect 12440 26367 12492 26376
rect 12440 26333 12449 26367
rect 12449 26333 12483 26367
rect 12483 26333 12492 26367
rect 12440 26324 12492 26333
rect 12716 26367 12768 26376
rect 12716 26333 12750 26367
rect 12750 26333 12768 26367
rect 12716 26324 12768 26333
rect 14096 26324 14148 26376
rect 17684 26392 17736 26444
rect 20536 26392 20588 26444
rect 4804 26256 4856 26308
rect 10508 26256 10560 26308
rect 14740 26256 14792 26308
rect 15568 26256 15620 26308
rect 18880 26324 18932 26376
rect 20904 26324 20956 26376
rect 21272 26367 21324 26376
rect 21272 26333 21281 26367
rect 21281 26333 21315 26367
rect 21315 26333 21324 26367
rect 21272 26324 21324 26333
rect 22100 26324 22152 26376
rect 3516 26188 3568 26240
rect 7104 26231 7156 26240
rect 7104 26197 7113 26231
rect 7113 26197 7147 26231
rect 7147 26197 7156 26231
rect 7104 26188 7156 26197
rect 9312 26231 9364 26240
rect 9312 26197 9321 26231
rect 9321 26197 9355 26231
rect 9355 26197 9364 26231
rect 9312 26188 9364 26197
rect 9404 26231 9456 26240
rect 9404 26197 9413 26231
rect 9413 26197 9447 26231
rect 9447 26197 9456 26231
rect 9404 26188 9456 26197
rect 13820 26231 13872 26240
rect 13820 26197 13829 26231
rect 13829 26197 13863 26231
rect 13863 26197 13872 26231
rect 13820 26188 13872 26197
rect 16120 26188 16172 26240
rect 16488 26256 16540 26308
rect 17960 26256 18012 26308
rect 19524 26299 19576 26308
rect 19524 26265 19533 26299
rect 19533 26265 19567 26299
rect 19567 26265 19576 26299
rect 19524 26256 19576 26265
rect 20260 26256 20312 26308
rect 23480 26256 23532 26308
rect 18052 26188 18104 26240
rect 21640 26188 21692 26240
rect 3658 26086 3710 26138
rect 3722 26086 3774 26138
rect 3786 26086 3838 26138
rect 3850 26086 3902 26138
rect 3914 26086 3966 26138
rect 3978 26086 4030 26138
rect 7658 26086 7710 26138
rect 7722 26086 7774 26138
rect 7786 26086 7838 26138
rect 7850 26086 7902 26138
rect 7914 26086 7966 26138
rect 7978 26086 8030 26138
rect 11658 26086 11710 26138
rect 11722 26086 11774 26138
rect 11786 26086 11838 26138
rect 11850 26086 11902 26138
rect 11914 26086 11966 26138
rect 11978 26086 12030 26138
rect 15658 26086 15710 26138
rect 15722 26086 15774 26138
rect 15786 26086 15838 26138
rect 15850 26086 15902 26138
rect 15914 26086 15966 26138
rect 15978 26086 16030 26138
rect 19658 26086 19710 26138
rect 19722 26086 19774 26138
rect 19786 26086 19838 26138
rect 19850 26086 19902 26138
rect 19914 26086 19966 26138
rect 19978 26086 20030 26138
rect 23658 26086 23710 26138
rect 23722 26086 23774 26138
rect 23786 26086 23838 26138
rect 23850 26086 23902 26138
rect 23914 26086 23966 26138
rect 23978 26086 24030 26138
rect 4988 25984 5040 26036
rect 9312 25984 9364 26036
rect 9772 25984 9824 26036
rect 10416 25984 10468 26036
rect 4436 25916 4488 25968
rect 6828 25916 6880 25968
rect 7104 25916 7156 25968
rect 11152 25916 11204 25968
rect 3516 25780 3568 25832
rect 5080 25848 5132 25900
rect 6092 25891 6144 25900
rect 6092 25857 6101 25891
rect 6101 25857 6135 25891
rect 6135 25857 6144 25891
rect 6092 25848 6144 25857
rect 7012 25891 7064 25900
rect 7012 25857 7021 25891
rect 7021 25857 7055 25891
rect 7055 25857 7064 25891
rect 7012 25848 7064 25857
rect 9036 25891 9088 25900
rect 9036 25857 9045 25891
rect 9045 25857 9079 25891
rect 9079 25857 9088 25891
rect 9036 25848 9088 25857
rect 4988 25780 5040 25832
rect 12256 25848 12308 25900
rect 15568 25984 15620 26036
rect 16672 25984 16724 26036
rect 17316 25984 17368 26036
rect 17684 25984 17736 26036
rect 13360 25916 13412 25968
rect 14648 25916 14700 25968
rect 15384 25916 15436 25968
rect 18052 26027 18104 26036
rect 18052 25993 18061 26027
rect 18061 25993 18095 26027
rect 18095 25993 18104 26027
rect 18052 25984 18104 25993
rect 18604 25984 18656 26036
rect 16120 25848 16172 25900
rect 17500 25891 17552 25900
rect 17500 25857 17509 25891
rect 17509 25857 17543 25891
rect 17543 25857 17552 25891
rect 17500 25848 17552 25857
rect 17684 25891 17736 25900
rect 17684 25857 17693 25891
rect 17693 25857 17727 25891
rect 17727 25857 17736 25891
rect 17684 25848 17736 25857
rect 18052 25848 18104 25900
rect 20076 25984 20128 26036
rect 22652 25984 22704 26036
rect 22100 25916 22152 25968
rect 23480 25916 23532 25968
rect 9680 25712 9732 25764
rect 9956 25712 10008 25764
rect 14280 25780 14332 25832
rect 17224 25823 17276 25832
rect 17224 25789 17233 25823
rect 17233 25789 17267 25823
rect 17267 25789 17276 25823
rect 17224 25780 17276 25789
rect 14464 25712 14516 25764
rect 16580 25712 16632 25764
rect 5172 25644 5224 25696
rect 5908 25687 5960 25696
rect 5908 25653 5917 25687
rect 5917 25653 5951 25687
rect 5951 25653 5960 25687
rect 5908 25644 5960 25653
rect 9220 25644 9272 25696
rect 10692 25644 10744 25696
rect 16304 25687 16356 25696
rect 16304 25653 16313 25687
rect 16313 25653 16347 25687
rect 16347 25653 16356 25687
rect 16304 25644 16356 25653
rect 16396 25644 16448 25696
rect 17868 25712 17920 25764
rect 18236 25712 18288 25764
rect 21364 25823 21416 25832
rect 21364 25789 21373 25823
rect 21373 25789 21407 25823
rect 21407 25789 21416 25823
rect 21364 25780 21416 25789
rect 22100 25780 22152 25832
rect 22468 25823 22520 25832
rect 22468 25789 22477 25823
rect 22477 25789 22511 25823
rect 22511 25789 22520 25823
rect 22468 25780 22520 25789
rect 23572 25712 23624 25764
rect 19340 25644 19392 25696
rect 2918 25542 2970 25594
rect 2982 25542 3034 25594
rect 3046 25542 3098 25594
rect 3110 25542 3162 25594
rect 3174 25542 3226 25594
rect 3238 25542 3290 25594
rect 6918 25542 6970 25594
rect 6982 25542 7034 25594
rect 7046 25542 7098 25594
rect 7110 25542 7162 25594
rect 7174 25542 7226 25594
rect 7238 25542 7290 25594
rect 10918 25542 10970 25594
rect 10982 25542 11034 25594
rect 11046 25542 11098 25594
rect 11110 25542 11162 25594
rect 11174 25542 11226 25594
rect 11238 25542 11290 25594
rect 14918 25542 14970 25594
rect 14982 25542 15034 25594
rect 15046 25542 15098 25594
rect 15110 25542 15162 25594
rect 15174 25542 15226 25594
rect 15238 25542 15290 25594
rect 18918 25542 18970 25594
rect 18982 25542 19034 25594
rect 19046 25542 19098 25594
rect 19110 25542 19162 25594
rect 19174 25542 19226 25594
rect 19238 25542 19290 25594
rect 22918 25542 22970 25594
rect 22982 25542 23034 25594
rect 23046 25542 23098 25594
rect 23110 25542 23162 25594
rect 23174 25542 23226 25594
rect 23238 25542 23290 25594
rect 4068 25483 4120 25492
rect 4068 25449 4077 25483
rect 4077 25449 4111 25483
rect 4111 25449 4120 25483
rect 4068 25440 4120 25449
rect 12992 25483 13044 25492
rect 12992 25449 13001 25483
rect 13001 25449 13035 25483
rect 13035 25449 13044 25483
rect 12992 25440 13044 25449
rect 15384 25440 15436 25492
rect 17960 25440 18012 25492
rect 19524 25440 19576 25492
rect 4988 25304 5040 25356
rect 7380 25347 7432 25356
rect 7380 25313 7389 25347
rect 7389 25313 7423 25347
rect 7423 25313 7432 25347
rect 7380 25304 7432 25313
rect 8852 25304 8904 25356
rect 12348 25304 12400 25356
rect 17868 25372 17920 25424
rect 22468 25372 22520 25424
rect 16488 25304 16540 25356
rect 18052 25304 18104 25356
rect 5448 25236 5500 25288
rect 5908 25236 5960 25288
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 9220 25236 9272 25288
rect 9956 25236 10008 25288
rect 5172 25168 5224 25220
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 13820 25236 13872 25288
rect 5908 25100 5960 25152
rect 6460 25100 6512 25152
rect 6552 25100 6604 25152
rect 10416 25168 10468 25220
rect 10508 25211 10560 25220
rect 10508 25177 10517 25211
rect 10517 25177 10551 25211
rect 10551 25177 10560 25211
rect 10508 25168 10560 25177
rect 10324 25100 10376 25152
rect 11520 25100 11572 25152
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 17408 25236 17460 25288
rect 18696 25236 18748 25288
rect 21180 25304 21232 25356
rect 21640 25347 21692 25356
rect 21640 25313 21649 25347
rect 21649 25313 21683 25347
rect 21683 25313 21692 25347
rect 21640 25304 21692 25313
rect 23572 25304 23624 25356
rect 16304 25168 16356 25220
rect 16212 25100 16264 25152
rect 17316 25100 17368 25152
rect 20536 25168 20588 25220
rect 20812 25211 20864 25220
rect 20812 25177 20821 25211
rect 20821 25177 20855 25211
rect 20855 25177 20864 25211
rect 20812 25168 20864 25177
rect 22560 25236 22612 25288
rect 20628 25100 20680 25152
rect 22652 25100 22704 25152
rect 3658 24998 3710 25050
rect 3722 24998 3774 25050
rect 3786 24998 3838 25050
rect 3850 24998 3902 25050
rect 3914 24998 3966 25050
rect 3978 24998 4030 25050
rect 7658 24998 7710 25050
rect 7722 24998 7774 25050
rect 7786 24998 7838 25050
rect 7850 24998 7902 25050
rect 7914 24998 7966 25050
rect 7978 24998 8030 25050
rect 11658 24998 11710 25050
rect 11722 24998 11774 25050
rect 11786 24998 11838 25050
rect 11850 24998 11902 25050
rect 11914 24998 11966 25050
rect 11978 24998 12030 25050
rect 15658 24998 15710 25050
rect 15722 24998 15774 25050
rect 15786 24998 15838 25050
rect 15850 24998 15902 25050
rect 15914 24998 15966 25050
rect 15978 24998 16030 25050
rect 19658 24998 19710 25050
rect 19722 24998 19774 25050
rect 19786 24998 19838 25050
rect 19850 24998 19902 25050
rect 19914 24998 19966 25050
rect 19978 24998 20030 25050
rect 23658 24998 23710 25050
rect 23722 24998 23774 25050
rect 23786 24998 23838 25050
rect 23850 24998 23902 25050
rect 23914 24998 23966 25050
rect 23978 24998 24030 25050
rect 6092 24896 6144 24948
rect 6460 24896 6512 24948
rect 6552 24828 6604 24880
rect 8852 24939 8904 24948
rect 8852 24905 8861 24939
rect 8861 24905 8895 24939
rect 8895 24905 8904 24939
rect 8852 24896 8904 24905
rect 9128 24896 9180 24948
rect 10508 24896 10560 24948
rect 15568 24896 15620 24948
rect 18052 24896 18104 24948
rect 9404 24828 9456 24880
rect 3516 24760 3568 24812
rect 5356 24760 5408 24812
rect 4988 24692 5040 24744
rect 4068 24624 4120 24676
rect 10324 24803 10376 24812
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 10508 24803 10560 24812
rect 10508 24769 10517 24803
rect 10517 24769 10551 24803
rect 10551 24769 10560 24803
rect 10508 24760 10560 24769
rect 7564 24692 7616 24744
rect 8668 24735 8720 24744
rect 8668 24701 8677 24735
rect 8677 24701 8711 24735
rect 8711 24701 8720 24735
rect 8668 24692 8720 24701
rect 8944 24692 8996 24744
rect 10692 24803 10744 24812
rect 10692 24769 10701 24803
rect 10701 24769 10735 24803
rect 10735 24769 10744 24803
rect 10692 24760 10744 24769
rect 13544 24760 13596 24812
rect 15568 24760 15620 24812
rect 19340 24760 19392 24812
rect 19524 24760 19576 24812
rect 11520 24692 11572 24744
rect 19892 24735 19944 24744
rect 19892 24701 19901 24735
rect 19901 24701 19935 24735
rect 19935 24701 19944 24735
rect 19892 24692 19944 24701
rect 21364 24692 21416 24744
rect 10324 24624 10376 24676
rect 10692 24624 10744 24676
rect 2136 24556 2188 24608
rect 3332 24556 3384 24608
rect 5264 24599 5316 24608
rect 5264 24565 5273 24599
rect 5273 24565 5307 24599
rect 5307 24565 5316 24599
rect 5264 24556 5316 24565
rect 19524 24556 19576 24608
rect 2918 24454 2970 24506
rect 2982 24454 3034 24506
rect 3046 24454 3098 24506
rect 3110 24454 3162 24506
rect 3174 24454 3226 24506
rect 3238 24454 3290 24506
rect 6918 24454 6970 24506
rect 6982 24454 7034 24506
rect 7046 24454 7098 24506
rect 7110 24454 7162 24506
rect 7174 24454 7226 24506
rect 7238 24454 7290 24506
rect 10918 24454 10970 24506
rect 10982 24454 11034 24506
rect 11046 24454 11098 24506
rect 11110 24454 11162 24506
rect 11174 24454 11226 24506
rect 11238 24454 11290 24506
rect 14918 24454 14970 24506
rect 14982 24454 15034 24506
rect 15046 24454 15098 24506
rect 15110 24454 15162 24506
rect 15174 24454 15226 24506
rect 15238 24454 15290 24506
rect 18918 24454 18970 24506
rect 18982 24454 19034 24506
rect 19046 24454 19098 24506
rect 19110 24454 19162 24506
rect 19174 24454 19226 24506
rect 19238 24454 19290 24506
rect 22918 24454 22970 24506
rect 22982 24454 23034 24506
rect 23046 24454 23098 24506
rect 23110 24454 23162 24506
rect 23174 24454 23226 24506
rect 23238 24454 23290 24506
rect 23480 24216 23532 24268
rect 1952 24148 2004 24200
rect 2136 24191 2188 24200
rect 2136 24157 2170 24191
rect 2170 24157 2188 24191
rect 2136 24148 2188 24157
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 4344 24080 4396 24132
rect 5448 24148 5500 24200
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 19892 24191 19944 24200
rect 19892 24157 19901 24191
rect 19901 24157 19935 24191
rect 19935 24157 19944 24191
rect 19892 24148 19944 24157
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 20168 24191 20220 24200
rect 20168 24157 20177 24191
rect 20177 24157 20211 24191
rect 20211 24157 20220 24191
rect 20168 24148 20220 24157
rect 22652 24148 22704 24200
rect 5264 24080 5316 24132
rect 7564 24080 7616 24132
rect 13544 24080 13596 24132
rect 3516 24012 3568 24064
rect 4620 24055 4672 24064
rect 4620 24021 4629 24055
rect 4629 24021 4663 24055
rect 4663 24021 4672 24055
rect 4620 24012 4672 24021
rect 6276 24055 6328 24064
rect 6276 24021 6285 24055
rect 6285 24021 6319 24055
rect 6319 24021 6328 24055
rect 6276 24012 6328 24021
rect 13176 24055 13228 24064
rect 13176 24021 13185 24055
rect 13185 24021 13219 24055
rect 13219 24021 13228 24055
rect 13176 24012 13228 24021
rect 22836 24080 22888 24132
rect 20260 24012 20312 24064
rect 21364 24012 21416 24064
rect 23204 24012 23256 24064
rect 25136 24080 25188 24132
rect 24492 24055 24544 24064
rect 24492 24021 24501 24055
rect 24501 24021 24535 24055
rect 24535 24021 24544 24055
rect 24492 24012 24544 24021
rect 3658 23910 3710 23962
rect 3722 23910 3774 23962
rect 3786 23910 3838 23962
rect 3850 23910 3902 23962
rect 3914 23910 3966 23962
rect 3978 23910 4030 23962
rect 7658 23910 7710 23962
rect 7722 23910 7774 23962
rect 7786 23910 7838 23962
rect 7850 23910 7902 23962
rect 7914 23910 7966 23962
rect 7978 23910 8030 23962
rect 11658 23910 11710 23962
rect 11722 23910 11774 23962
rect 11786 23910 11838 23962
rect 11850 23910 11902 23962
rect 11914 23910 11966 23962
rect 11978 23910 12030 23962
rect 15658 23910 15710 23962
rect 15722 23910 15774 23962
rect 15786 23910 15838 23962
rect 15850 23910 15902 23962
rect 15914 23910 15966 23962
rect 15978 23910 16030 23962
rect 19658 23910 19710 23962
rect 19722 23910 19774 23962
rect 19786 23910 19838 23962
rect 19850 23910 19902 23962
rect 19914 23910 19966 23962
rect 19978 23910 20030 23962
rect 23658 23910 23710 23962
rect 23722 23910 23774 23962
rect 23786 23910 23838 23962
rect 23850 23910 23902 23962
rect 23914 23910 23966 23962
rect 23978 23910 24030 23962
rect 4068 23808 4120 23860
rect 4804 23808 4856 23860
rect 6828 23851 6880 23860
rect 6828 23817 6837 23851
rect 6837 23817 6871 23851
rect 6871 23817 6880 23851
rect 6828 23808 6880 23817
rect 4620 23783 4672 23792
rect 1952 23672 2004 23724
rect 4620 23749 4654 23783
rect 4654 23749 4672 23783
rect 4620 23740 4672 23749
rect 4988 23740 5040 23792
rect 12808 23740 12860 23792
rect 13452 23808 13504 23860
rect 20076 23808 20128 23860
rect 4068 23672 4120 23724
rect 4344 23715 4396 23724
rect 4344 23681 4353 23715
rect 4353 23681 4387 23715
rect 4387 23681 4396 23715
rect 4344 23672 4396 23681
rect 5724 23579 5776 23588
rect 5724 23545 5733 23579
rect 5733 23545 5767 23579
rect 5767 23545 5776 23579
rect 7380 23672 7432 23724
rect 12256 23672 12308 23724
rect 7472 23604 7524 23656
rect 7564 23604 7616 23656
rect 5724 23536 5776 23545
rect 6828 23536 6880 23588
rect 8116 23604 8168 23656
rect 8392 23604 8444 23656
rect 12440 23604 12492 23656
rect 12808 23579 12860 23588
rect 12808 23545 12817 23579
rect 12817 23545 12851 23579
rect 12851 23545 12860 23579
rect 12808 23536 12860 23545
rect 6000 23468 6052 23520
rect 8760 23468 8812 23520
rect 11336 23468 11388 23520
rect 14280 23511 14332 23520
rect 14280 23477 14289 23511
rect 14289 23477 14323 23511
rect 14323 23477 14332 23511
rect 16948 23740 17000 23792
rect 17224 23740 17276 23792
rect 17960 23740 18012 23792
rect 19248 23740 19300 23792
rect 19708 23740 19760 23792
rect 15568 23604 15620 23656
rect 16672 23715 16724 23724
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 18420 23672 18472 23724
rect 18328 23604 18380 23656
rect 14280 23468 14332 23477
rect 16764 23468 16816 23520
rect 18420 23468 18472 23520
rect 18512 23468 18564 23520
rect 19432 23468 19484 23520
rect 19892 23715 19944 23724
rect 19892 23681 19901 23715
rect 19901 23681 19935 23715
rect 19935 23681 19944 23715
rect 22100 23740 22152 23792
rect 19892 23672 19944 23681
rect 20536 23672 20588 23724
rect 20260 23604 20312 23656
rect 22376 23647 22428 23656
rect 22376 23613 22385 23647
rect 22385 23613 22419 23647
rect 22419 23613 22428 23647
rect 22376 23604 22428 23613
rect 22836 23647 22888 23656
rect 22836 23613 22845 23647
rect 22845 23613 22879 23647
rect 22879 23613 22888 23647
rect 22836 23604 22888 23613
rect 20904 23536 20956 23588
rect 23204 23715 23256 23724
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 24492 23740 24544 23792
rect 23388 23604 23440 23656
rect 19800 23468 19852 23520
rect 23572 23468 23624 23520
rect 25136 23468 25188 23520
rect 2918 23366 2970 23418
rect 2982 23366 3034 23418
rect 3046 23366 3098 23418
rect 3110 23366 3162 23418
rect 3174 23366 3226 23418
rect 3238 23366 3290 23418
rect 6918 23366 6970 23418
rect 6982 23366 7034 23418
rect 7046 23366 7098 23418
rect 7110 23366 7162 23418
rect 7174 23366 7226 23418
rect 7238 23366 7290 23418
rect 10918 23366 10970 23418
rect 10982 23366 11034 23418
rect 11046 23366 11098 23418
rect 11110 23366 11162 23418
rect 11174 23366 11226 23418
rect 11238 23366 11290 23418
rect 14918 23366 14970 23418
rect 14982 23366 15034 23418
rect 15046 23366 15098 23418
rect 15110 23366 15162 23418
rect 15174 23366 15226 23418
rect 15238 23366 15290 23418
rect 18918 23366 18970 23418
rect 18982 23366 19034 23418
rect 19046 23366 19098 23418
rect 19110 23366 19162 23418
rect 19174 23366 19226 23418
rect 19238 23366 19290 23418
rect 22918 23366 22970 23418
rect 22982 23366 23034 23418
rect 23046 23366 23098 23418
rect 23110 23366 23162 23418
rect 23174 23366 23226 23418
rect 23238 23366 23290 23418
rect 5356 23264 5408 23316
rect 7380 23264 7432 23316
rect 5540 23196 5592 23248
rect 10876 23264 10928 23316
rect 12164 23307 12216 23316
rect 12164 23273 12173 23307
rect 12173 23273 12207 23307
rect 12207 23273 12216 23307
rect 12164 23264 12216 23273
rect 12256 23264 12308 23316
rect 8576 23196 8628 23248
rect 1952 23171 2004 23180
rect 1952 23137 1961 23171
rect 1961 23137 1995 23171
rect 1995 23137 2004 23171
rect 1952 23128 2004 23137
rect 5724 23128 5776 23180
rect 5908 23171 5960 23180
rect 5908 23137 5917 23171
rect 5917 23137 5951 23171
rect 5951 23137 5960 23171
rect 5908 23128 5960 23137
rect 6000 23171 6052 23180
rect 6000 23137 6009 23171
rect 6009 23137 6043 23171
rect 6043 23137 6052 23171
rect 6000 23128 6052 23137
rect 7380 23128 7432 23180
rect 5080 23103 5132 23112
rect 5080 23069 5089 23103
rect 5089 23069 5123 23103
rect 5123 23069 5132 23103
rect 5080 23060 5132 23069
rect 5448 23060 5500 23112
rect 6276 23103 6328 23112
rect 6276 23069 6285 23103
rect 6285 23069 6319 23103
rect 6319 23069 6328 23103
rect 6276 23060 6328 23069
rect 6552 23103 6604 23112
rect 6552 23069 6561 23103
rect 6561 23069 6595 23103
rect 6595 23069 6604 23103
rect 6552 23060 6604 23069
rect 9680 23128 9732 23180
rect 10416 23171 10468 23180
rect 10416 23137 10425 23171
rect 10425 23137 10459 23171
rect 10459 23137 10468 23171
rect 10416 23128 10468 23137
rect 12256 23128 12308 23180
rect 8668 23060 8720 23112
rect 8760 23103 8812 23112
rect 8760 23069 8769 23103
rect 8769 23069 8803 23103
rect 8803 23069 8812 23103
rect 8760 23060 8812 23069
rect 9496 23060 9548 23112
rect 10324 23060 10376 23112
rect 14832 23264 14884 23316
rect 17316 23264 17368 23316
rect 12440 23196 12492 23248
rect 16672 23171 16724 23180
rect 16672 23137 16681 23171
rect 16681 23137 16715 23171
rect 16715 23137 16724 23171
rect 16672 23128 16724 23137
rect 18420 23128 18472 23180
rect 13176 23060 13228 23112
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 15568 23060 15620 23112
rect 16120 23103 16172 23112
rect 16120 23069 16127 23103
rect 16127 23069 16172 23103
rect 16120 23060 16172 23069
rect 16304 23103 16356 23112
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 17408 23060 17460 23112
rect 18328 23060 18380 23112
rect 19892 23264 19944 23316
rect 21732 23264 21784 23316
rect 19524 23196 19576 23248
rect 19984 23196 20036 23248
rect 22376 23196 22428 23248
rect 20536 23128 20588 23180
rect 22100 23128 22152 23180
rect 22744 23128 22796 23180
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 19800 23103 19852 23112
rect 19800 23069 19809 23103
rect 19809 23069 19843 23103
rect 19843 23069 19852 23103
rect 19800 23060 19852 23069
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 2320 22992 2372 23044
rect 5264 22992 5316 23044
rect 7380 22992 7432 23044
rect 7564 22992 7616 23044
rect 3148 22924 3200 22976
rect 5356 22967 5408 22976
rect 5356 22933 5365 22967
rect 5365 22933 5399 22967
rect 5399 22933 5408 22967
rect 5356 22924 5408 22933
rect 6184 22924 6236 22976
rect 10140 22924 10192 22976
rect 10324 22967 10376 22976
rect 10324 22933 10333 22967
rect 10333 22933 10367 22967
rect 10367 22933 10376 22967
rect 10324 22924 10376 22933
rect 10692 23035 10744 23044
rect 10692 23001 10701 23035
rect 10701 23001 10735 23035
rect 10735 23001 10744 23035
rect 10692 22992 10744 23001
rect 12900 22992 12952 23044
rect 11428 22924 11480 22976
rect 13728 22924 13780 22976
rect 14372 23035 14424 23044
rect 14372 23001 14406 23035
rect 14406 23001 14424 23035
rect 14372 22992 14424 23001
rect 18052 22992 18104 23044
rect 18420 23035 18472 23044
rect 18420 23001 18429 23035
rect 18429 23001 18463 23035
rect 18463 23001 18472 23035
rect 18420 22992 18472 23001
rect 18972 22992 19024 23044
rect 20812 23103 20864 23112
rect 20812 23069 20821 23103
rect 20821 23069 20855 23103
rect 20855 23069 20864 23103
rect 20812 23060 20864 23069
rect 20904 23060 20956 23112
rect 22192 23103 22244 23112
rect 22192 23069 22201 23103
rect 22201 23069 22235 23103
rect 22235 23069 22244 23103
rect 22192 23060 22244 23069
rect 21088 22992 21140 23044
rect 15476 22967 15528 22976
rect 15476 22933 15485 22967
rect 15485 22933 15519 22967
rect 15519 22933 15528 22967
rect 15476 22924 15528 22933
rect 16120 22924 16172 22976
rect 16488 22924 16540 22976
rect 16580 22967 16632 22976
rect 16580 22933 16589 22967
rect 16589 22933 16623 22967
rect 16623 22933 16632 22967
rect 16580 22924 16632 22933
rect 19432 22924 19484 22976
rect 20352 22967 20404 22976
rect 20352 22933 20379 22967
rect 20379 22933 20404 22967
rect 20352 22924 20404 22933
rect 20996 22967 21048 22976
rect 20996 22933 21005 22967
rect 21005 22933 21039 22967
rect 21039 22933 21048 22967
rect 20996 22924 21048 22933
rect 24216 22967 24268 22976
rect 24216 22933 24225 22967
rect 24225 22933 24259 22967
rect 24259 22933 24268 22967
rect 24216 22924 24268 22933
rect 24492 22967 24544 22976
rect 24492 22933 24501 22967
rect 24501 22933 24535 22967
rect 24535 22933 24544 22967
rect 24492 22924 24544 22933
rect 3658 22822 3710 22874
rect 3722 22822 3774 22874
rect 3786 22822 3838 22874
rect 3850 22822 3902 22874
rect 3914 22822 3966 22874
rect 3978 22822 4030 22874
rect 7658 22822 7710 22874
rect 7722 22822 7774 22874
rect 7786 22822 7838 22874
rect 7850 22822 7902 22874
rect 7914 22822 7966 22874
rect 7978 22822 8030 22874
rect 11658 22822 11710 22874
rect 11722 22822 11774 22874
rect 11786 22822 11838 22874
rect 11850 22822 11902 22874
rect 11914 22822 11966 22874
rect 11978 22822 12030 22874
rect 15658 22822 15710 22874
rect 15722 22822 15774 22874
rect 15786 22822 15838 22874
rect 15850 22822 15902 22874
rect 15914 22822 15966 22874
rect 15978 22822 16030 22874
rect 19658 22822 19710 22874
rect 19722 22822 19774 22874
rect 19786 22822 19838 22874
rect 19850 22822 19902 22874
rect 19914 22822 19966 22874
rect 19978 22822 20030 22874
rect 23658 22822 23710 22874
rect 23722 22822 23774 22874
rect 23786 22822 23838 22874
rect 23850 22822 23902 22874
rect 23914 22822 23966 22874
rect 23978 22822 24030 22874
rect 2320 22763 2372 22772
rect 2320 22729 2329 22763
rect 2329 22729 2363 22763
rect 2363 22729 2372 22763
rect 2320 22720 2372 22729
rect 3148 22763 3200 22772
rect 3148 22729 3157 22763
rect 3157 22729 3191 22763
rect 3191 22729 3200 22763
rect 3148 22720 3200 22729
rect 3332 22652 3384 22704
rect 3516 22584 3568 22636
rect 4620 22652 4672 22704
rect 9496 22763 9548 22772
rect 9496 22729 9505 22763
rect 9505 22729 9539 22763
rect 9539 22729 9548 22763
rect 9496 22720 9548 22729
rect 10692 22720 10744 22772
rect 8300 22695 8352 22704
rect 8300 22661 8309 22695
rect 8309 22661 8343 22695
rect 8343 22661 8352 22695
rect 8300 22652 8352 22661
rect 8576 22652 8628 22704
rect 11336 22652 11388 22704
rect 12164 22720 12216 22772
rect 13360 22763 13412 22772
rect 13360 22729 13369 22763
rect 13369 22729 13403 22763
rect 13403 22729 13412 22763
rect 13360 22720 13412 22729
rect 13728 22763 13780 22772
rect 13728 22729 13737 22763
rect 13737 22729 13771 22763
rect 13771 22729 13780 22763
rect 13728 22720 13780 22729
rect 14372 22763 14424 22772
rect 14372 22729 14381 22763
rect 14381 22729 14415 22763
rect 14415 22729 14424 22763
rect 14372 22720 14424 22729
rect 12256 22652 12308 22704
rect 3976 22627 4028 22636
rect 3976 22593 3985 22627
rect 3985 22593 4019 22627
rect 4019 22593 4028 22627
rect 3976 22584 4028 22593
rect 7380 22584 7432 22636
rect 7472 22584 7524 22636
rect 4436 22516 4488 22568
rect 6460 22516 6512 22568
rect 8760 22584 8812 22636
rect 9588 22627 9640 22636
rect 9588 22593 9597 22627
rect 9597 22593 9631 22627
rect 9631 22593 9640 22627
rect 9588 22584 9640 22593
rect 9496 22516 9548 22568
rect 10324 22516 10376 22568
rect 10416 22516 10468 22568
rect 11980 22584 12032 22636
rect 11428 22516 11480 22568
rect 4528 22380 4580 22432
rect 8024 22423 8076 22432
rect 8024 22389 8033 22423
rect 8033 22389 8067 22423
rect 8067 22389 8076 22423
rect 8024 22380 8076 22389
rect 8852 22380 8904 22432
rect 9128 22423 9180 22432
rect 9128 22389 9137 22423
rect 9137 22389 9171 22423
rect 9171 22389 9180 22423
rect 9128 22380 9180 22389
rect 9956 22380 10008 22432
rect 12624 22559 12676 22568
rect 12624 22525 12633 22559
rect 12633 22525 12667 22559
rect 12667 22525 12676 22559
rect 12624 22516 12676 22525
rect 12900 22695 12952 22704
rect 12900 22661 12909 22695
rect 12909 22661 12943 22695
rect 12943 22661 12952 22695
rect 12900 22652 12952 22661
rect 13452 22584 13504 22636
rect 13636 22584 13688 22636
rect 15476 22720 15528 22772
rect 16212 22652 16264 22704
rect 16672 22695 16724 22704
rect 16672 22661 16681 22695
rect 16681 22661 16715 22695
rect 16715 22661 16724 22695
rect 16672 22652 16724 22661
rect 17960 22652 18012 22704
rect 18972 22652 19024 22704
rect 19432 22695 19484 22704
rect 19432 22661 19441 22695
rect 19441 22661 19475 22695
rect 19475 22661 19484 22695
rect 19432 22652 19484 22661
rect 13544 22516 13596 22568
rect 16120 22584 16172 22636
rect 17316 22584 17368 22636
rect 20168 22720 20220 22772
rect 22192 22720 22244 22772
rect 20076 22652 20128 22704
rect 14280 22448 14332 22500
rect 14832 22448 14884 22500
rect 12716 22380 12768 22432
rect 13728 22380 13780 22432
rect 17684 22559 17736 22568
rect 17684 22525 17693 22559
rect 17693 22525 17727 22559
rect 17727 22525 17736 22559
rect 17684 22516 17736 22525
rect 20168 22584 20220 22636
rect 24216 22652 24268 22704
rect 24492 22652 24544 22704
rect 20444 22584 20496 22636
rect 21088 22584 21140 22636
rect 21732 22584 21784 22636
rect 23388 22584 23440 22636
rect 25228 22584 25280 22636
rect 20720 22516 20772 22568
rect 21548 22516 21600 22568
rect 20352 22380 20404 22432
rect 20536 22448 20588 22500
rect 21180 22448 21232 22500
rect 21916 22448 21968 22500
rect 22284 22559 22336 22568
rect 22284 22525 22293 22559
rect 22293 22525 22327 22559
rect 22327 22525 22336 22559
rect 22284 22516 22336 22525
rect 23940 22559 23992 22568
rect 23940 22525 23949 22559
rect 23949 22525 23983 22559
rect 23983 22525 23992 22559
rect 23940 22516 23992 22525
rect 23480 22448 23532 22500
rect 26516 22491 26568 22500
rect 26516 22457 26525 22491
rect 26525 22457 26559 22491
rect 26559 22457 26568 22491
rect 26516 22448 26568 22457
rect 25412 22423 25464 22432
rect 25412 22389 25421 22423
rect 25421 22389 25455 22423
rect 25455 22389 25464 22423
rect 25412 22380 25464 22389
rect 2918 22278 2970 22330
rect 2982 22278 3034 22330
rect 3046 22278 3098 22330
rect 3110 22278 3162 22330
rect 3174 22278 3226 22330
rect 3238 22278 3290 22330
rect 6918 22278 6970 22330
rect 6982 22278 7034 22330
rect 7046 22278 7098 22330
rect 7110 22278 7162 22330
rect 7174 22278 7226 22330
rect 7238 22278 7290 22330
rect 10918 22278 10970 22330
rect 10982 22278 11034 22330
rect 11046 22278 11098 22330
rect 11110 22278 11162 22330
rect 11174 22278 11226 22330
rect 11238 22278 11290 22330
rect 14918 22278 14970 22330
rect 14982 22278 15034 22330
rect 15046 22278 15098 22330
rect 15110 22278 15162 22330
rect 15174 22278 15226 22330
rect 15238 22278 15290 22330
rect 18918 22278 18970 22330
rect 18982 22278 19034 22330
rect 19046 22278 19098 22330
rect 19110 22278 19162 22330
rect 19174 22278 19226 22330
rect 19238 22278 19290 22330
rect 22918 22278 22970 22330
rect 22982 22278 23034 22330
rect 23046 22278 23098 22330
rect 23110 22278 23162 22330
rect 23174 22278 23226 22330
rect 23238 22278 23290 22330
rect 7380 22176 7432 22228
rect 9128 22176 9180 22228
rect 3976 22108 4028 22160
rect 4252 22108 4304 22160
rect 8760 22108 8812 22160
rect 12624 22176 12676 22228
rect 15568 22176 15620 22228
rect 17868 22176 17920 22228
rect 19524 22176 19576 22228
rect 20076 22176 20128 22228
rect 12716 22108 12768 22160
rect 13912 22108 13964 22160
rect 4344 22040 4396 22092
rect 6460 22040 6512 22092
rect 8208 22040 8260 22092
rect 8668 22040 8720 22092
rect 2688 22015 2740 22024
rect 2688 21981 2697 22015
rect 2697 21981 2731 22015
rect 2731 21981 2740 22015
rect 2688 21972 2740 21981
rect 4896 22015 4948 22024
rect 4896 21981 4905 22015
rect 4905 21981 4939 22015
rect 4939 21981 4948 22015
rect 4896 21972 4948 21981
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 4620 21904 4672 21956
rect 8024 21972 8076 22024
rect 8576 22015 8628 22024
rect 8576 21981 8585 22015
rect 8585 21981 8619 22015
rect 8619 21981 8628 22015
rect 8576 21972 8628 21981
rect 15476 22040 15528 22092
rect 17316 22040 17368 22092
rect 12440 21972 12492 22024
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 5448 21904 5500 21956
rect 2320 21836 2372 21888
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 5908 21836 5960 21888
rect 8116 21836 8168 21888
rect 11152 21904 11204 21956
rect 15384 21947 15436 21956
rect 15384 21913 15393 21947
rect 15393 21913 15427 21947
rect 15427 21913 15436 21947
rect 15384 21904 15436 21913
rect 15476 21947 15528 21956
rect 15476 21913 15485 21947
rect 15485 21913 15519 21947
rect 15519 21913 15528 21947
rect 15476 21904 15528 21913
rect 16764 21972 16816 22024
rect 18512 22015 18564 22024
rect 17132 21904 17184 21956
rect 18512 21981 18521 22015
rect 18521 21981 18555 22015
rect 18555 21981 18564 22015
rect 18512 21972 18564 21981
rect 17592 21904 17644 21956
rect 17868 21904 17920 21956
rect 18328 21904 18380 21956
rect 19248 22040 19300 22092
rect 18696 21972 18748 22024
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 9496 21836 9548 21888
rect 17684 21836 17736 21888
rect 20076 21972 20128 22024
rect 22284 22176 22336 22228
rect 23940 22176 23992 22228
rect 20904 22108 20956 22160
rect 21916 22151 21968 22160
rect 21916 22117 21925 22151
rect 21925 22117 21959 22151
rect 21959 22117 21968 22151
rect 21916 22108 21968 22117
rect 23480 22108 23532 22160
rect 25228 22040 25280 22092
rect 19524 21836 19576 21888
rect 21548 22015 21600 22024
rect 21548 21981 21557 22015
rect 21557 21981 21591 22015
rect 21591 21981 21600 22015
rect 21548 21972 21600 21981
rect 21732 22015 21784 22024
rect 21732 21981 21741 22015
rect 21741 21981 21775 22015
rect 21775 21981 21784 22015
rect 21732 21972 21784 21981
rect 22192 22015 22244 22024
rect 22192 21981 22201 22015
rect 22201 21981 22235 22015
rect 22235 21981 22244 22015
rect 22192 21972 22244 21981
rect 24124 21904 24176 21956
rect 20812 21879 20864 21888
rect 20812 21845 20821 21879
rect 20821 21845 20855 21879
rect 20855 21845 20864 21879
rect 20812 21836 20864 21845
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 24400 22015 24452 22024
rect 24400 21981 24409 22015
rect 24409 21981 24443 22015
rect 24443 21981 24452 22015
rect 24400 21972 24452 21981
rect 3658 21734 3710 21786
rect 3722 21734 3774 21786
rect 3786 21734 3838 21786
rect 3850 21734 3902 21786
rect 3914 21734 3966 21786
rect 3978 21734 4030 21786
rect 7658 21734 7710 21786
rect 7722 21734 7774 21786
rect 7786 21734 7838 21786
rect 7850 21734 7902 21786
rect 7914 21734 7966 21786
rect 7978 21734 8030 21786
rect 11658 21734 11710 21786
rect 11722 21734 11774 21786
rect 11786 21734 11838 21786
rect 11850 21734 11902 21786
rect 11914 21734 11966 21786
rect 11978 21734 12030 21786
rect 15658 21734 15710 21786
rect 15722 21734 15774 21786
rect 15786 21734 15838 21786
rect 15850 21734 15902 21786
rect 15914 21734 15966 21786
rect 15978 21734 16030 21786
rect 19658 21734 19710 21786
rect 19722 21734 19774 21786
rect 19786 21734 19838 21786
rect 19850 21734 19902 21786
rect 19914 21734 19966 21786
rect 19978 21734 20030 21786
rect 23658 21734 23710 21786
rect 23722 21734 23774 21786
rect 23786 21734 23838 21786
rect 23850 21734 23902 21786
rect 23914 21734 23966 21786
rect 23978 21734 24030 21786
rect 1952 21496 2004 21548
rect 2320 21539 2372 21548
rect 2320 21505 2354 21539
rect 2354 21505 2372 21539
rect 2320 21496 2372 21505
rect 4712 21564 4764 21616
rect 5356 21564 5408 21616
rect 8576 21632 8628 21684
rect 9496 21675 9548 21684
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 4344 21496 4396 21548
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 8208 21564 8260 21616
rect 10048 21564 10100 21616
rect 6368 21539 6420 21548
rect 6368 21505 6377 21539
rect 6377 21505 6411 21539
rect 6411 21505 6420 21539
rect 6368 21496 6420 21505
rect 6000 21471 6052 21480
rect 6000 21437 6009 21471
rect 6009 21437 6043 21471
rect 6043 21437 6052 21471
rect 6000 21428 6052 21437
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 6828 21539 6880 21548
rect 6828 21505 6842 21539
rect 6842 21505 6876 21539
rect 6876 21505 6880 21539
rect 6828 21496 6880 21505
rect 8944 21496 8996 21548
rect 9404 21428 9456 21480
rect 12624 21632 12676 21684
rect 15476 21632 15528 21684
rect 17960 21632 18012 21684
rect 19248 21632 19300 21684
rect 19616 21632 19668 21684
rect 21272 21675 21324 21684
rect 21272 21641 21281 21675
rect 21281 21641 21315 21675
rect 21315 21641 21324 21675
rect 21272 21632 21324 21641
rect 21732 21632 21784 21684
rect 24400 21632 24452 21684
rect 20536 21564 20588 21616
rect 12256 21496 12308 21548
rect 14096 21496 14148 21548
rect 14464 21539 14516 21548
rect 14464 21505 14498 21539
rect 14498 21505 14516 21539
rect 14464 21496 14516 21505
rect 16304 21496 16356 21548
rect 12348 21428 12400 21480
rect 16212 21471 16264 21480
rect 16212 21437 16221 21471
rect 16221 21437 16255 21471
rect 16255 21437 16264 21471
rect 16212 21428 16264 21437
rect 18604 21428 18656 21480
rect 20352 21539 20404 21548
rect 20352 21505 20361 21539
rect 20361 21505 20395 21539
rect 20395 21505 20404 21539
rect 22192 21564 22244 21616
rect 20352 21496 20404 21505
rect 21180 21539 21232 21548
rect 21180 21505 21189 21539
rect 21189 21505 21223 21539
rect 21223 21505 21232 21539
rect 21180 21496 21232 21505
rect 22652 21496 22704 21548
rect 24768 21496 24820 21548
rect 18420 21360 18472 21412
rect 20260 21360 20312 21412
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 23480 21428 23532 21480
rect 24124 21428 24176 21480
rect 24584 21428 24636 21480
rect 25412 21496 25464 21548
rect 26056 21496 26108 21548
rect 21364 21360 21416 21412
rect 3516 21292 3568 21344
rect 3976 21292 4028 21344
rect 5632 21335 5684 21344
rect 5632 21301 5641 21335
rect 5641 21301 5675 21335
rect 5675 21301 5684 21335
rect 5632 21292 5684 21301
rect 5724 21335 5776 21344
rect 5724 21301 5733 21335
rect 5733 21301 5767 21335
rect 5767 21301 5776 21335
rect 5724 21292 5776 21301
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 6644 21292 6696 21344
rect 15568 21292 15620 21344
rect 15660 21335 15712 21344
rect 15660 21301 15669 21335
rect 15669 21301 15703 21335
rect 15703 21301 15712 21335
rect 15660 21292 15712 21301
rect 20168 21292 20220 21344
rect 20812 21292 20864 21344
rect 21916 21335 21968 21344
rect 21916 21301 21925 21335
rect 21925 21301 21959 21335
rect 21959 21301 21968 21335
rect 21916 21292 21968 21301
rect 24216 21292 24268 21344
rect 24952 21292 25004 21344
rect 25504 21292 25556 21344
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 2918 21190 2970 21242
rect 2982 21190 3034 21242
rect 3046 21190 3098 21242
rect 3110 21190 3162 21242
rect 3174 21190 3226 21242
rect 3238 21190 3290 21242
rect 6918 21190 6970 21242
rect 6982 21190 7034 21242
rect 7046 21190 7098 21242
rect 7110 21190 7162 21242
rect 7174 21190 7226 21242
rect 7238 21190 7290 21242
rect 10918 21190 10970 21242
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 11238 21190 11290 21242
rect 14918 21190 14970 21242
rect 14982 21190 15034 21242
rect 15046 21190 15098 21242
rect 15110 21190 15162 21242
rect 15174 21190 15226 21242
rect 15238 21190 15290 21242
rect 18918 21190 18970 21242
rect 18982 21190 19034 21242
rect 19046 21190 19098 21242
rect 19110 21190 19162 21242
rect 19174 21190 19226 21242
rect 19238 21190 19290 21242
rect 22918 21190 22970 21242
rect 22982 21190 23034 21242
rect 23046 21190 23098 21242
rect 23110 21190 23162 21242
rect 23174 21190 23226 21242
rect 23238 21190 23290 21242
rect 2688 21088 2740 21140
rect 4436 21088 4488 21140
rect 8208 21088 8260 21140
rect 10232 21088 10284 21140
rect 14464 21088 14516 21140
rect 1952 20995 2004 21004
rect 1952 20961 1961 20995
rect 1961 20961 1995 20995
rect 1995 20961 2004 20995
rect 1952 20952 2004 20961
rect 6460 20995 6512 21004
rect 6460 20961 6469 20995
rect 6469 20961 6503 20995
rect 6503 20961 6512 20995
rect 6460 20952 6512 20961
rect 19616 21088 19668 21140
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 18512 21020 18564 21072
rect 3976 20884 4028 20936
rect 5724 20884 5776 20936
rect 9588 20927 9640 20936
rect 9588 20893 9597 20927
rect 9597 20893 9631 20927
rect 9631 20893 9640 20927
rect 9588 20884 9640 20893
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 15660 20884 15712 20936
rect 16948 20927 17000 20936
rect 16948 20893 16957 20927
rect 16957 20893 16991 20927
rect 16991 20893 17000 20927
rect 16948 20884 17000 20893
rect 17132 20927 17184 20936
rect 17132 20893 17141 20927
rect 17141 20893 17175 20927
rect 17175 20893 17184 20927
rect 17132 20884 17184 20893
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 18328 20927 18380 20936
rect 18328 20893 18337 20927
rect 18337 20893 18371 20927
rect 18371 20893 18380 20927
rect 18328 20884 18380 20893
rect 18604 20927 18656 20936
rect 18604 20893 18613 20927
rect 18613 20893 18647 20927
rect 18647 20893 18656 20927
rect 18604 20884 18656 20893
rect 19432 20952 19484 21004
rect 22100 21020 22152 21072
rect 2412 20816 2464 20868
rect 5540 20816 5592 20868
rect 6736 20859 6788 20868
rect 6736 20825 6770 20859
rect 6770 20825 6788 20859
rect 6736 20816 6788 20825
rect 18144 20816 18196 20868
rect 18788 20816 18840 20868
rect 19524 20816 19576 20868
rect 20260 20927 20312 20936
rect 20260 20893 20269 20927
rect 20269 20893 20303 20927
rect 20303 20893 20312 20927
rect 20260 20884 20312 20893
rect 3332 20791 3384 20800
rect 3332 20757 3341 20791
rect 3341 20757 3375 20791
rect 3375 20757 3384 20791
rect 3332 20748 3384 20757
rect 4160 20748 4212 20800
rect 5816 20748 5868 20800
rect 7380 20748 7432 20800
rect 8760 20748 8812 20800
rect 15568 20748 15620 20800
rect 18696 20748 18748 20800
rect 20444 20748 20496 20800
rect 23480 20884 23532 20936
rect 24768 20884 24820 20936
rect 22192 20791 22244 20800
rect 22192 20757 22201 20791
rect 22201 20757 22235 20791
rect 22235 20757 22244 20791
rect 22192 20748 22244 20757
rect 23572 20748 23624 20800
rect 24216 20816 24268 20868
rect 25688 20816 25740 20868
rect 26148 20816 26200 20868
rect 24124 20791 24176 20800
rect 24124 20757 24133 20791
rect 24133 20757 24167 20791
rect 24167 20757 24176 20791
rect 24124 20748 24176 20757
rect 3658 20646 3710 20698
rect 3722 20646 3774 20698
rect 3786 20646 3838 20698
rect 3850 20646 3902 20698
rect 3914 20646 3966 20698
rect 3978 20646 4030 20698
rect 7658 20646 7710 20698
rect 7722 20646 7774 20698
rect 7786 20646 7838 20698
rect 7850 20646 7902 20698
rect 7914 20646 7966 20698
rect 7978 20646 8030 20698
rect 11658 20646 11710 20698
rect 11722 20646 11774 20698
rect 11786 20646 11838 20698
rect 11850 20646 11902 20698
rect 11914 20646 11966 20698
rect 11978 20646 12030 20698
rect 15658 20646 15710 20698
rect 15722 20646 15774 20698
rect 15786 20646 15838 20698
rect 15850 20646 15902 20698
rect 15914 20646 15966 20698
rect 15978 20646 16030 20698
rect 19658 20646 19710 20698
rect 19722 20646 19774 20698
rect 19786 20646 19838 20698
rect 19850 20646 19902 20698
rect 19914 20646 19966 20698
rect 19978 20646 20030 20698
rect 23658 20646 23710 20698
rect 23722 20646 23774 20698
rect 23786 20646 23838 20698
rect 23850 20646 23902 20698
rect 23914 20646 23966 20698
rect 23978 20646 24030 20698
rect 2412 20587 2464 20596
rect 2412 20553 2421 20587
rect 2421 20553 2455 20587
rect 2455 20553 2464 20587
rect 2412 20544 2464 20553
rect 3332 20544 3384 20596
rect 4896 20587 4948 20596
rect 4896 20553 4905 20587
rect 4905 20553 4939 20587
rect 4939 20553 4948 20587
rect 4896 20544 4948 20553
rect 5632 20544 5684 20596
rect 6736 20587 6788 20596
rect 6736 20553 6745 20587
rect 6745 20553 6779 20587
rect 6779 20553 6788 20587
rect 6736 20544 6788 20553
rect 3516 20476 3568 20528
rect 5816 20476 5868 20528
rect 3976 20451 4028 20460
rect 3976 20417 3985 20451
rect 3985 20417 4019 20451
rect 4019 20417 4028 20451
rect 3976 20408 4028 20417
rect 4252 20408 4304 20460
rect 5264 20408 5316 20460
rect 3516 20383 3568 20392
rect 3516 20349 3525 20383
rect 3525 20349 3559 20383
rect 3559 20349 3568 20383
rect 3516 20340 3568 20349
rect 7380 20587 7432 20596
rect 7380 20553 7389 20587
rect 7389 20553 7423 20587
rect 7423 20553 7432 20587
rect 7380 20544 7432 20553
rect 7656 20544 7708 20596
rect 12808 20544 12860 20596
rect 15384 20544 15436 20596
rect 8208 20476 8260 20528
rect 12256 20476 12308 20528
rect 10324 20408 10376 20460
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 13728 20408 13780 20460
rect 14004 20451 14056 20460
rect 14004 20417 14011 20451
rect 14011 20417 14056 20451
rect 14004 20408 14056 20417
rect 10048 20340 10100 20392
rect 13452 20340 13504 20392
rect 4160 20272 4212 20324
rect 6368 20272 6420 20324
rect 16488 20476 16540 20528
rect 18604 20544 18656 20596
rect 18328 20476 18380 20528
rect 20260 20544 20312 20596
rect 19524 20476 19576 20528
rect 19616 20476 19668 20528
rect 14372 20408 14424 20460
rect 3976 20204 4028 20256
rect 14280 20272 14332 20324
rect 8576 20204 8628 20256
rect 13084 20247 13136 20256
rect 13084 20213 13093 20247
rect 13093 20213 13127 20247
rect 13127 20213 13136 20247
rect 13084 20204 13136 20213
rect 13360 20247 13412 20256
rect 13360 20213 13369 20247
rect 13369 20213 13403 20247
rect 13403 20213 13412 20247
rect 13360 20204 13412 20213
rect 13912 20204 13964 20256
rect 18512 20408 18564 20460
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 19340 20408 19392 20460
rect 19892 20451 19944 20460
rect 19892 20417 19901 20451
rect 19901 20417 19935 20451
rect 19935 20417 19944 20451
rect 19892 20408 19944 20417
rect 20168 20408 20220 20460
rect 20444 20519 20496 20528
rect 20444 20485 20453 20519
rect 20453 20485 20487 20519
rect 20487 20485 20496 20519
rect 20444 20476 20496 20485
rect 20720 20408 20772 20460
rect 22652 20451 22704 20460
rect 22652 20417 22661 20451
rect 22661 20417 22695 20451
rect 22695 20417 22704 20451
rect 22652 20408 22704 20417
rect 24400 20544 24452 20596
rect 24952 20544 25004 20596
rect 24124 20519 24176 20528
rect 24124 20485 24133 20519
rect 24133 20485 24167 20519
rect 24167 20485 24176 20519
rect 24124 20476 24176 20485
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 17868 20383 17920 20392
rect 17868 20349 17877 20383
rect 17877 20349 17911 20383
rect 17911 20349 17920 20383
rect 17868 20340 17920 20349
rect 18144 20340 18196 20392
rect 18328 20383 18380 20392
rect 18328 20349 18337 20383
rect 18337 20349 18371 20383
rect 18371 20349 18380 20383
rect 18328 20340 18380 20349
rect 18420 20340 18472 20392
rect 19708 20340 19760 20392
rect 19800 20340 19852 20392
rect 20352 20340 20404 20392
rect 20904 20383 20956 20392
rect 20904 20349 20913 20383
rect 20913 20349 20947 20383
rect 20947 20349 20956 20383
rect 20904 20340 20956 20349
rect 22192 20340 22244 20392
rect 22560 20340 22612 20392
rect 25504 20451 25556 20460
rect 25504 20417 25513 20451
rect 25513 20417 25547 20451
rect 25547 20417 25556 20451
rect 25504 20408 25556 20417
rect 25780 20408 25832 20460
rect 24124 20340 24176 20392
rect 24676 20340 24728 20392
rect 26424 20340 26476 20392
rect 18788 20204 18840 20256
rect 19524 20204 19576 20256
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 22008 20247 22060 20256
rect 22008 20213 22017 20247
rect 22017 20213 22051 20247
rect 22051 20213 22060 20247
rect 22008 20204 22060 20213
rect 23480 20204 23532 20256
rect 23664 20247 23716 20256
rect 23664 20213 23673 20247
rect 23673 20213 23707 20247
rect 23707 20213 23716 20247
rect 23664 20204 23716 20213
rect 24400 20247 24452 20256
rect 24400 20213 24409 20247
rect 24409 20213 24443 20247
rect 24443 20213 24452 20247
rect 24400 20204 24452 20213
rect 25228 20204 25280 20256
rect 2918 20102 2970 20154
rect 2982 20102 3034 20154
rect 3046 20102 3098 20154
rect 3110 20102 3162 20154
rect 3174 20102 3226 20154
rect 3238 20102 3290 20154
rect 6918 20102 6970 20154
rect 6982 20102 7034 20154
rect 7046 20102 7098 20154
rect 7110 20102 7162 20154
rect 7174 20102 7226 20154
rect 7238 20102 7290 20154
rect 10918 20102 10970 20154
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 11238 20102 11290 20154
rect 14918 20102 14970 20154
rect 14982 20102 15034 20154
rect 15046 20102 15098 20154
rect 15110 20102 15162 20154
rect 15174 20102 15226 20154
rect 15238 20102 15290 20154
rect 18918 20102 18970 20154
rect 18982 20102 19034 20154
rect 19046 20102 19098 20154
rect 19110 20102 19162 20154
rect 19174 20102 19226 20154
rect 19238 20102 19290 20154
rect 22918 20102 22970 20154
rect 22982 20102 23034 20154
rect 23046 20102 23098 20154
rect 23110 20102 23162 20154
rect 23174 20102 23226 20154
rect 23238 20102 23290 20154
rect 2504 19796 2556 19848
rect 3148 19796 3200 19848
rect 3976 19839 4028 19848
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 5172 20000 5224 20052
rect 7012 20000 7064 20052
rect 7656 20000 7708 20052
rect 13268 20000 13320 20052
rect 13728 19932 13780 19984
rect 20260 20000 20312 20052
rect 8668 19864 8720 19916
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 6644 19796 6696 19848
rect 8576 19839 8628 19848
rect 8576 19805 8585 19839
rect 8585 19805 8619 19839
rect 8619 19805 8628 19839
rect 8576 19796 8628 19805
rect 14188 19864 14240 19916
rect 10968 19796 11020 19848
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 13360 19796 13412 19848
rect 14004 19796 14056 19848
rect 16948 19864 17000 19916
rect 16764 19796 16816 19848
rect 18144 19864 18196 19916
rect 18972 19864 19024 19916
rect 19616 19864 19668 19916
rect 19708 19864 19760 19916
rect 20352 19864 20404 19916
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22008 19864 22060 19873
rect 22468 19907 22520 19916
rect 22468 19873 22477 19907
rect 22477 19873 22511 19907
rect 22511 19873 22520 19907
rect 22468 19864 22520 19873
rect 17592 19796 17644 19848
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 2412 19728 2464 19780
rect 6552 19728 6604 19780
rect 4804 19660 4856 19712
rect 6092 19660 6144 19712
rect 6736 19660 6788 19712
rect 7196 19660 7248 19712
rect 8116 19703 8168 19712
rect 8116 19669 8125 19703
rect 8125 19669 8159 19703
rect 8159 19669 8168 19703
rect 8116 19660 8168 19669
rect 11520 19728 11572 19780
rect 13636 19728 13688 19780
rect 14648 19728 14700 19780
rect 18328 19728 18380 19780
rect 18420 19728 18472 19780
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 19800 19839 19852 19848
rect 19800 19805 19809 19839
rect 19809 19805 19843 19839
rect 19843 19805 19852 19839
rect 19800 19796 19852 19805
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 23572 20000 23624 20052
rect 24676 20043 24728 20052
rect 24676 20009 24685 20043
rect 24685 20009 24719 20043
rect 24719 20009 24728 20043
rect 24676 20000 24728 20009
rect 24400 19932 24452 19984
rect 25504 19932 25556 19984
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 12164 19660 12216 19712
rect 13360 19660 13412 19712
rect 14280 19660 14332 19712
rect 16488 19660 16540 19712
rect 17592 19660 17644 19712
rect 19340 19728 19392 19780
rect 20444 19728 20496 19780
rect 21916 19728 21968 19780
rect 22100 19728 22152 19780
rect 24124 19796 24176 19848
rect 25228 19839 25280 19848
rect 25228 19805 25237 19839
rect 25237 19805 25271 19839
rect 25271 19805 25280 19839
rect 25228 19796 25280 19805
rect 25780 19796 25832 19848
rect 20260 19660 20312 19712
rect 26424 19660 26476 19712
rect 3658 19558 3710 19610
rect 3722 19558 3774 19610
rect 3786 19558 3838 19610
rect 3850 19558 3902 19610
rect 3914 19558 3966 19610
rect 3978 19558 4030 19610
rect 7658 19558 7710 19610
rect 7722 19558 7774 19610
rect 7786 19558 7838 19610
rect 7850 19558 7902 19610
rect 7914 19558 7966 19610
rect 7978 19558 8030 19610
rect 11658 19558 11710 19610
rect 11722 19558 11774 19610
rect 11786 19558 11838 19610
rect 11850 19558 11902 19610
rect 11914 19558 11966 19610
rect 11978 19558 12030 19610
rect 15658 19558 15710 19610
rect 15722 19558 15774 19610
rect 15786 19558 15838 19610
rect 15850 19558 15902 19610
rect 15914 19558 15966 19610
rect 15978 19558 16030 19610
rect 19658 19558 19710 19610
rect 19722 19558 19774 19610
rect 19786 19558 19838 19610
rect 19850 19558 19902 19610
rect 19914 19558 19966 19610
rect 19978 19558 20030 19610
rect 23658 19558 23710 19610
rect 23722 19558 23774 19610
rect 23786 19558 23838 19610
rect 23850 19558 23902 19610
rect 23914 19558 23966 19610
rect 23978 19558 24030 19610
rect 2412 19499 2464 19508
rect 2412 19465 2421 19499
rect 2421 19465 2455 19499
rect 2455 19465 2464 19499
rect 2412 19456 2464 19465
rect 3148 19499 3200 19508
rect 3148 19465 3157 19499
rect 3157 19465 3191 19499
rect 3191 19465 3200 19499
rect 3148 19456 3200 19465
rect 6552 19499 6604 19508
rect 6552 19465 6561 19499
rect 6561 19465 6595 19499
rect 6595 19465 6604 19499
rect 6552 19456 6604 19465
rect 4068 19388 4120 19440
rect 4712 19431 4764 19440
rect 4712 19397 4721 19431
rect 4721 19397 4755 19431
rect 4755 19397 4764 19431
rect 4712 19388 4764 19397
rect 6460 19388 6512 19440
rect 3332 19320 3384 19372
rect 4252 19320 4304 19372
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 8116 19456 8168 19508
rect 10324 19456 10376 19508
rect 7012 19431 7064 19440
rect 7012 19397 7021 19431
rect 7021 19397 7055 19431
rect 7055 19397 7064 19431
rect 7012 19388 7064 19397
rect 7104 19431 7156 19440
rect 7104 19397 7113 19431
rect 7113 19397 7147 19431
rect 7147 19397 7156 19431
rect 7104 19388 7156 19397
rect 7380 19388 7432 19440
rect 3516 19252 3568 19304
rect 7196 19363 7248 19372
rect 7196 19329 7210 19363
rect 7210 19329 7244 19363
rect 7244 19329 7248 19363
rect 7196 19320 7248 19329
rect 8208 19320 8260 19372
rect 7380 19227 7432 19236
rect 7380 19193 7389 19227
rect 7389 19193 7423 19227
rect 7423 19193 7432 19227
rect 7380 19184 7432 19193
rect 8116 19295 8168 19304
rect 8116 19261 8125 19295
rect 8125 19261 8159 19295
rect 8159 19261 8168 19295
rect 8116 19252 8168 19261
rect 8760 19388 8812 19440
rect 10968 19388 11020 19440
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 12256 19499 12308 19508
rect 12256 19465 12265 19499
rect 12265 19465 12299 19499
rect 12299 19465 12308 19499
rect 12256 19456 12308 19465
rect 13544 19456 13596 19508
rect 14280 19456 14332 19508
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 18052 19456 18104 19508
rect 20168 19456 20220 19508
rect 21180 19456 21232 19508
rect 22468 19456 22520 19508
rect 13084 19388 13136 19440
rect 14096 19388 14148 19440
rect 9956 19363 10008 19372
rect 9956 19329 9965 19363
rect 9965 19329 9999 19363
rect 9999 19329 10008 19363
rect 9956 19320 10008 19329
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 7564 19184 7616 19236
rect 9680 19184 9732 19236
rect 10232 19295 10284 19304
rect 10232 19261 10241 19295
rect 10241 19261 10275 19295
rect 10275 19261 10284 19295
rect 10232 19252 10284 19261
rect 10692 19252 10744 19304
rect 11428 19184 11480 19236
rect 11888 19320 11940 19372
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 12532 19320 12584 19372
rect 14004 19320 14056 19372
rect 16764 19431 16816 19440
rect 16764 19397 16773 19431
rect 16773 19397 16807 19431
rect 16807 19397 16816 19431
rect 16764 19388 16816 19397
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 9128 19159 9180 19168
rect 9128 19125 9137 19159
rect 9137 19125 9171 19159
rect 9171 19125 9180 19159
rect 9128 19116 9180 19125
rect 9312 19116 9364 19168
rect 16948 19320 17000 19372
rect 18420 19388 18472 19440
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 18604 19320 18656 19372
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19524 19363 19576 19372
rect 19524 19329 19533 19363
rect 19533 19329 19567 19363
rect 19567 19329 19576 19363
rect 19524 19320 19576 19329
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 20076 19320 20128 19372
rect 20352 19320 20404 19372
rect 22192 19320 22244 19372
rect 14280 19116 14332 19168
rect 20168 19252 20220 19304
rect 22652 19252 22704 19304
rect 19524 19116 19576 19168
rect 22100 19116 22152 19168
rect 2918 19014 2970 19066
rect 2982 19014 3034 19066
rect 3046 19014 3098 19066
rect 3110 19014 3162 19066
rect 3174 19014 3226 19066
rect 3238 19014 3290 19066
rect 6918 19014 6970 19066
rect 6982 19014 7034 19066
rect 7046 19014 7098 19066
rect 7110 19014 7162 19066
rect 7174 19014 7226 19066
rect 7238 19014 7290 19066
rect 10918 19014 10970 19066
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 11238 19014 11290 19066
rect 14918 19014 14970 19066
rect 14982 19014 15034 19066
rect 15046 19014 15098 19066
rect 15110 19014 15162 19066
rect 15174 19014 15226 19066
rect 15238 19014 15290 19066
rect 18918 19014 18970 19066
rect 18982 19014 19034 19066
rect 19046 19014 19098 19066
rect 19110 19014 19162 19066
rect 19174 19014 19226 19066
rect 19238 19014 19290 19066
rect 22918 19014 22970 19066
rect 22982 19014 23034 19066
rect 23046 19014 23098 19066
rect 23110 19014 23162 19066
rect 23174 19014 23226 19066
rect 23238 19014 23290 19066
rect 4988 18912 5040 18964
rect 9128 18912 9180 18964
rect 9864 18912 9916 18964
rect 9956 18912 10008 18964
rect 10784 18912 10836 18964
rect 12072 18912 12124 18964
rect 5080 18776 5132 18828
rect 6552 18776 6604 18828
rect 3516 18708 3568 18760
rect 2136 18615 2188 18624
rect 2136 18581 2145 18615
rect 2145 18581 2179 18615
rect 2179 18581 2188 18615
rect 2136 18572 2188 18581
rect 2780 18572 2832 18624
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 4896 18751 4948 18760
rect 4896 18717 4906 18751
rect 4906 18717 4940 18751
rect 4940 18717 4948 18751
rect 4896 18708 4948 18717
rect 5264 18751 5316 18760
rect 5264 18717 5278 18751
rect 5278 18717 5312 18751
rect 5312 18717 5316 18751
rect 5264 18708 5316 18717
rect 7196 18708 7248 18760
rect 7472 18708 7524 18760
rect 10692 18844 10744 18896
rect 17040 18912 17092 18964
rect 22192 18955 22244 18964
rect 22192 18921 22201 18955
rect 22201 18921 22235 18955
rect 22235 18921 22244 18955
rect 22192 18912 22244 18921
rect 26424 18955 26476 18964
rect 26424 18921 26433 18955
rect 26433 18921 26467 18955
rect 26467 18921 26476 18955
rect 26424 18912 26476 18921
rect 8760 18776 8812 18828
rect 4344 18683 4396 18692
rect 4344 18649 4353 18683
rect 4353 18649 4387 18683
rect 4387 18649 4396 18683
rect 4344 18640 4396 18649
rect 4252 18572 4304 18624
rect 4988 18640 5040 18692
rect 7564 18640 7616 18692
rect 8484 18708 8536 18760
rect 9312 18708 9364 18760
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 14096 18776 14148 18828
rect 8208 18683 8260 18692
rect 8208 18649 8217 18683
rect 8217 18649 8251 18683
rect 8251 18649 8260 18683
rect 8208 18640 8260 18649
rect 9128 18640 9180 18692
rect 5540 18572 5592 18624
rect 6920 18572 6972 18624
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 8300 18572 8352 18624
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 12072 18708 12124 18760
rect 14372 18708 14424 18760
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 18144 18776 18196 18828
rect 19340 18776 19392 18828
rect 18604 18708 18656 18760
rect 22560 18708 22612 18760
rect 23388 18708 23440 18760
rect 12992 18640 13044 18692
rect 15108 18640 15160 18692
rect 17500 18640 17552 18692
rect 17684 18683 17736 18692
rect 17684 18649 17693 18683
rect 17693 18649 17727 18683
rect 17727 18649 17736 18683
rect 17684 18640 17736 18649
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 16856 18572 16908 18624
rect 18696 18640 18748 18692
rect 18880 18640 18932 18692
rect 25044 18640 25096 18692
rect 26240 18640 26292 18692
rect 19708 18572 19760 18624
rect 3658 18470 3710 18522
rect 3722 18470 3774 18522
rect 3786 18470 3838 18522
rect 3850 18470 3902 18522
rect 3914 18470 3966 18522
rect 3978 18470 4030 18522
rect 7658 18470 7710 18522
rect 7722 18470 7774 18522
rect 7786 18470 7838 18522
rect 7850 18470 7902 18522
rect 7914 18470 7966 18522
rect 7978 18470 8030 18522
rect 11658 18470 11710 18522
rect 11722 18470 11774 18522
rect 11786 18470 11838 18522
rect 11850 18470 11902 18522
rect 11914 18470 11966 18522
rect 11978 18470 12030 18522
rect 15658 18470 15710 18522
rect 15722 18470 15774 18522
rect 15786 18470 15838 18522
rect 15850 18470 15902 18522
rect 15914 18470 15966 18522
rect 15978 18470 16030 18522
rect 19658 18470 19710 18522
rect 19722 18470 19774 18522
rect 19786 18470 19838 18522
rect 19850 18470 19902 18522
rect 19914 18470 19966 18522
rect 19978 18470 20030 18522
rect 23658 18470 23710 18522
rect 23722 18470 23774 18522
rect 23786 18470 23838 18522
rect 23850 18470 23902 18522
rect 23914 18470 23966 18522
rect 23978 18470 24030 18522
rect 4344 18368 4396 18420
rect 5356 18411 5408 18420
rect 5356 18377 5365 18411
rect 5365 18377 5399 18411
rect 5399 18377 5408 18411
rect 5356 18368 5408 18377
rect 2504 18275 2556 18284
rect 2504 18241 2513 18275
rect 2513 18241 2547 18275
rect 2547 18241 2556 18275
rect 2504 18232 2556 18241
rect 2780 18275 2832 18284
rect 2780 18241 2814 18275
rect 2814 18241 2832 18275
rect 2780 18232 2832 18241
rect 4068 18232 4120 18284
rect 5632 18275 5684 18284
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 7012 18368 7064 18420
rect 7472 18368 7524 18420
rect 8300 18368 8352 18420
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 7104 18232 7156 18284
rect 8024 18232 8076 18284
rect 8208 18232 8260 18284
rect 9211 18343 9263 18352
rect 9211 18309 9220 18343
rect 9220 18309 9254 18343
rect 9254 18309 9263 18343
rect 9211 18300 9263 18309
rect 9772 18368 9824 18420
rect 15108 18411 15160 18420
rect 15108 18377 15117 18411
rect 15117 18377 15151 18411
rect 15151 18377 15160 18411
rect 15108 18368 15160 18377
rect 9680 18300 9732 18352
rect 8576 18207 8628 18216
rect 8576 18173 8585 18207
rect 8585 18173 8619 18207
rect 8619 18173 8628 18207
rect 8576 18164 8628 18173
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 12072 18164 12124 18216
rect 14740 18164 14792 18216
rect 16396 18300 16448 18352
rect 18144 18300 18196 18352
rect 18880 18343 18932 18352
rect 18880 18309 18889 18343
rect 18889 18309 18923 18343
rect 18923 18309 18932 18343
rect 18880 18300 18932 18309
rect 16856 18232 16908 18284
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 16396 18207 16448 18216
rect 16396 18173 16405 18207
rect 16405 18173 16439 18207
rect 16439 18173 16448 18207
rect 16396 18164 16448 18173
rect 16764 18207 16816 18216
rect 16764 18173 16773 18207
rect 16773 18173 16807 18207
rect 16807 18173 16816 18207
rect 16764 18164 16816 18173
rect 18420 18275 18472 18284
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 22100 18232 22152 18284
rect 23388 18368 23440 18420
rect 23848 18300 23900 18352
rect 25780 18411 25832 18420
rect 25780 18377 25789 18411
rect 25789 18377 25823 18411
rect 25823 18377 25832 18411
rect 25780 18368 25832 18377
rect 26240 18411 26292 18420
rect 26240 18377 26249 18411
rect 26249 18377 26283 18411
rect 26283 18377 26292 18411
rect 26240 18368 26292 18377
rect 24860 18300 24912 18352
rect 26056 18275 26108 18284
rect 26056 18241 26065 18275
rect 26065 18241 26099 18275
rect 26099 18241 26108 18275
rect 26056 18232 26108 18241
rect 18604 18164 18656 18216
rect 4160 18028 4212 18080
rect 5172 18028 5224 18080
rect 7104 18028 7156 18080
rect 7196 18028 7248 18080
rect 8116 18028 8168 18080
rect 14832 18096 14884 18148
rect 16120 18096 16172 18148
rect 17040 18096 17092 18148
rect 17776 18096 17828 18148
rect 18144 18096 18196 18148
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 23480 18164 23532 18216
rect 9956 18028 10008 18080
rect 15384 18028 15436 18080
rect 17868 18028 17920 18080
rect 24124 18028 24176 18080
rect 25964 18071 26016 18080
rect 25964 18037 25973 18071
rect 25973 18037 26007 18071
rect 26007 18037 26016 18071
rect 25964 18028 26016 18037
rect 2918 17926 2970 17978
rect 2982 17926 3034 17978
rect 3046 17926 3098 17978
rect 3110 17926 3162 17978
rect 3174 17926 3226 17978
rect 3238 17926 3290 17978
rect 6918 17926 6970 17978
rect 6982 17926 7034 17978
rect 7046 17926 7098 17978
rect 7110 17926 7162 17978
rect 7174 17926 7226 17978
rect 7238 17926 7290 17978
rect 10918 17926 10970 17978
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 11238 17926 11290 17978
rect 14918 17926 14970 17978
rect 14982 17926 15034 17978
rect 15046 17926 15098 17978
rect 15110 17926 15162 17978
rect 15174 17926 15226 17978
rect 15238 17926 15290 17978
rect 18918 17926 18970 17978
rect 18982 17926 19034 17978
rect 19046 17926 19098 17978
rect 19110 17926 19162 17978
rect 19174 17926 19226 17978
rect 19238 17926 19290 17978
rect 22918 17926 22970 17978
rect 22982 17926 23034 17978
rect 23046 17926 23098 17978
rect 23110 17926 23162 17978
rect 23174 17926 23226 17978
rect 23238 17926 23290 17978
rect 3516 17824 3568 17876
rect 5632 17824 5684 17876
rect 8024 17867 8076 17876
rect 8024 17833 8033 17867
rect 8033 17833 8067 17867
rect 8067 17833 8076 17867
rect 8024 17824 8076 17833
rect 8576 17824 8628 17876
rect 9220 17824 9272 17876
rect 9496 17824 9548 17876
rect 10324 17824 10376 17876
rect 10600 17824 10652 17876
rect 17224 17824 17276 17876
rect 17684 17824 17736 17876
rect 1492 17663 1544 17672
rect 1492 17629 1501 17663
rect 1501 17629 1535 17663
rect 1535 17629 1544 17663
rect 1492 17620 1544 17629
rect 2136 17620 2188 17672
rect 6552 17756 6604 17808
rect 11428 17756 11480 17808
rect 4344 17731 4396 17740
rect 4344 17697 4353 17731
rect 4353 17697 4387 17731
rect 4387 17697 4396 17731
rect 4344 17688 4396 17697
rect 4896 17620 4948 17672
rect 5356 17620 5408 17672
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 5448 17552 5500 17604
rect 6644 17731 6696 17740
rect 6644 17697 6653 17731
rect 6653 17697 6687 17731
rect 6687 17697 6696 17731
rect 6644 17688 6696 17697
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 10784 17688 10836 17740
rect 12256 17688 12308 17740
rect 14004 17688 14056 17740
rect 18604 17731 18656 17740
rect 18604 17697 18613 17731
rect 18613 17697 18647 17731
rect 18647 17697 18656 17731
rect 18604 17688 18656 17697
rect 22100 17824 22152 17876
rect 23480 17824 23532 17876
rect 23848 17867 23900 17876
rect 23848 17833 23857 17867
rect 23857 17833 23891 17867
rect 23891 17833 23900 17867
rect 23848 17824 23900 17833
rect 24860 17824 24912 17876
rect 26148 17867 26200 17876
rect 26148 17833 26157 17867
rect 26157 17833 26191 17867
rect 26191 17833 26200 17867
rect 26148 17824 26200 17833
rect 22284 17688 22336 17740
rect 22560 17688 22612 17740
rect 6920 17663 6972 17672
rect 6920 17629 6954 17663
rect 6954 17629 6972 17663
rect 6920 17620 6972 17629
rect 9772 17663 9824 17672
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 13176 17620 13228 17672
rect 14372 17620 14424 17672
rect 16764 17620 16816 17672
rect 8944 17552 8996 17604
rect 10692 17595 10744 17604
rect 10692 17561 10701 17595
rect 10701 17561 10735 17595
rect 10735 17561 10744 17595
rect 10692 17552 10744 17561
rect 17960 17620 18012 17672
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 23388 17688 23440 17740
rect 19340 17552 19392 17604
rect 4804 17484 4856 17536
rect 9772 17484 9824 17536
rect 11336 17484 11388 17536
rect 12808 17484 12860 17536
rect 16120 17484 16172 17536
rect 17500 17484 17552 17536
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 26056 17620 26108 17672
rect 24768 17552 24820 17604
rect 26056 17484 26108 17536
rect 3658 17382 3710 17434
rect 3722 17382 3774 17434
rect 3786 17382 3838 17434
rect 3850 17382 3902 17434
rect 3914 17382 3966 17434
rect 3978 17382 4030 17434
rect 7658 17382 7710 17434
rect 7722 17382 7774 17434
rect 7786 17382 7838 17434
rect 7850 17382 7902 17434
rect 7914 17382 7966 17434
rect 7978 17382 8030 17434
rect 11658 17382 11710 17434
rect 11722 17382 11774 17434
rect 11786 17382 11838 17434
rect 11850 17382 11902 17434
rect 11914 17382 11966 17434
rect 11978 17382 12030 17434
rect 15658 17382 15710 17434
rect 15722 17382 15774 17434
rect 15786 17382 15838 17434
rect 15850 17382 15902 17434
rect 15914 17382 15966 17434
rect 15978 17382 16030 17434
rect 19658 17382 19710 17434
rect 19722 17382 19774 17434
rect 19786 17382 19838 17434
rect 19850 17382 19902 17434
rect 19914 17382 19966 17434
rect 19978 17382 20030 17434
rect 23658 17382 23710 17434
rect 23722 17382 23774 17434
rect 23786 17382 23838 17434
rect 23850 17382 23902 17434
rect 23914 17382 23966 17434
rect 23978 17382 24030 17434
rect 1492 17212 1544 17264
rect 2504 17212 2556 17264
rect 12992 17323 13044 17332
rect 12992 17289 13001 17323
rect 13001 17289 13035 17323
rect 13035 17289 13044 17323
rect 12992 17280 13044 17289
rect 4620 17212 4672 17264
rect 6736 17212 6788 17264
rect 10232 17212 10284 17264
rect 2228 17144 2280 17196
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4804 17144 4856 17196
rect 9680 17144 9732 17196
rect 10508 17187 10560 17196
rect 10508 17153 10517 17187
rect 10517 17153 10551 17187
rect 10551 17153 10560 17187
rect 10508 17144 10560 17153
rect 2780 17008 2832 17060
rect 3516 17008 3568 17060
rect 4344 17076 4396 17128
rect 12624 17119 12676 17128
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 8944 17008 8996 17060
rect 9496 17008 9548 17060
rect 12900 17076 12952 17128
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 17132 17212 17184 17264
rect 19340 17280 19392 17332
rect 22468 17280 22520 17332
rect 25044 17280 25096 17332
rect 19432 17212 19484 17264
rect 22836 17212 22888 17264
rect 23388 17212 23440 17264
rect 25964 17212 26016 17264
rect 13728 17144 13780 17196
rect 14372 17144 14424 17196
rect 14556 17187 14608 17196
rect 14556 17153 14590 17187
rect 14590 17153 14608 17187
rect 14556 17144 14608 17153
rect 13820 17076 13872 17128
rect 4436 16940 4488 16992
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 11520 16940 11572 16992
rect 15476 16940 15528 16992
rect 16028 17187 16080 17196
rect 16028 17153 16037 17187
rect 16037 17153 16071 17187
rect 16071 17153 16080 17187
rect 16028 17144 16080 17153
rect 16120 17187 16172 17196
rect 16120 17153 16129 17187
rect 16129 17153 16163 17187
rect 16163 17153 16172 17187
rect 16120 17144 16172 17153
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 16488 17076 16540 17128
rect 16764 17076 16816 17128
rect 17684 17076 17736 17128
rect 21548 17076 21600 17128
rect 22560 17076 22612 17128
rect 26056 17119 26108 17128
rect 26056 17085 26065 17119
rect 26065 17085 26099 17119
rect 26099 17085 26108 17119
rect 26056 17076 26108 17085
rect 16672 16940 16724 16992
rect 19432 16940 19484 16992
rect 21456 16940 21508 16992
rect 22100 16940 22152 16992
rect 2918 16838 2970 16890
rect 2982 16838 3034 16890
rect 3046 16838 3098 16890
rect 3110 16838 3162 16890
rect 3174 16838 3226 16890
rect 3238 16838 3290 16890
rect 6918 16838 6970 16890
rect 6982 16838 7034 16890
rect 7046 16838 7098 16890
rect 7110 16838 7162 16890
rect 7174 16838 7226 16890
rect 7238 16838 7290 16890
rect 10918 16838 10970 16890
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 11238 16838 11290 16890
rect 14918 16838 14970 16890
rect 14982 16838 15034 16890
rect 15046 16838 15098 16890
rect 15110 16838 15162 16890
rect 15174 16838 15226 16890
rect 15238 16838 15290 16890
rect 18918 16838 18970 16890
rect 18982 16838 19034 16890
rect 19046 16838 19098 16890
rect 19110 16838 19162 16890
rect 19174 16838 19226 16890
rect 19238 16838 19290 16890
rect 22918 16838 22970 16890
rect 22982 16838 23034 16890
rect 23046 16838 23098 16890
rect 23110 16838 23162 16890
rect 23174 16838 23226 16890
rect 23238 16838 23290 16890
rect 2228 16779 2280 16788
rect 2228 16745 2237 16779
rect 2237 16745 2271 16779
rect 2271 16745 2280 16779
rect 2228 16736 2280 16745
rect 6000 16736 6052 16788
rect 9680 16736 9732 16788
rect 4988 16600 5040 16652
rect 8208 16668 8260 16720
rect 10692 16736 10744 16788
rect 13268 16736 13320 16788
rect 13820 16779 13872 16788
rect 13820 16745 13829 16779
rect 13829 16745 13863 16779
rect 13863 16745 13872 16779
rect 13820 16736 13872 16745
rect 10968 16668 11020 16720
rect 16488 16736 16540 16788
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 2780 16532 2832 16584
rect 4252 16575 4304 16584
rect 4252 16541 4261 16575
rect 4261 16541 4295 16575
rect 4295 16541 4304 16575
rect 4252 16532 4304 16541
rect 4344 16575 4396 16584
rect 4344 16541 4354 16575
rect 4354 16541 4388 16575
rect 4388 16541 4396 16575
rect 4344 16532 4396 16541
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 5356 16532 5408 16584
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 4988 16464 5040 16516
rect 7288 16507 7340 16516
rect 7288 16473 7297 16507
rect 7297 16473 7331 16507
rect 7331 16473 7340 16507
rect 7288 16464 7340 16473
rect 7380 16507 7432 16516
rect 7380 16473 7389 16507
rect 7389 16473 7423 16507
rect 7423 16473 7432 16507
rect 7380 16464 7432 16473
rect 10324 16532 10376 16584
rect 11336 16532 11388 16584
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 13176 16532 13228 16584
rect 14832 16600 14884 16652
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 5264 16396 5316 16448
rect 5908 16396 5960 16448
rect 7564 16396 7616 16448
rect 11428 16439 11480 16448
rect 11428 16405 11437 16439
rect 11437 16405 11471 16439
rect 11471 16405 11480 16439
rect 11428 16396 11480 16405
rect 12256 16464 12308 16516
rect 13544 16507 13596 16516
rect 13544 16473 13553 16507
rect 13553 16473 13587 16507
rect 13587 16473 13596 16507
rect 13544 16464 13596 16473
rect 14372 16532 14424 16584
rect 16580 16600 16632 16652
rect 18420 16736 18472 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 20076 16779 20128 16788
rect 20076 16745 20085 16779
rect 20085 16745 20119 16779
rect 20119 16745 20128 16779
rect 20076 16736 20128 16745
rect 19616 16668 19668 16720
rect 14280 16396 14332 16448
rect 16028 16532 16080 16584
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 18696 16600 18748 16652
rect 20628 16668 20680 16720
rect 22100 16736 22152 16788
rect 17592 16532 17644 16584
rect 18788 16532 18840 16584
rect 19248 16532 19300 16584
rect 19432 16532 19484 16584
rect 20996 16643 21048 16652
rect 20996 16609 21005 16643
rect 21005 16609 21039 16643
rect 21039 16609 21048 16643
rect 20996 16600 21048 16609
rect 21548 16600 21600 16652
rect 20352 16575 20404 16584
rect 20352 16541 20361 16575
rect 20361 16541 20395 16575
rect 20395 16541 20404 16575
rect 20352 16532 20404 16541
rect 15568 16507 15620 16516
rect 15568 16473 15602 16507
rect 15602 16473 15620 16507
rect 15568 16464 15620 16473
rect 14740 16396 14792 16448
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 17040 16464 17092 16516
rect 17960 16507 18012 16516
rect 17960 16473 17994 16507
rect 17994 16473 18012 16507
rect 17960 16464 18012 16473
rect 16764 16439 16816 16448
rect 16764 16405 16773 16439
rect 16773 16405 16807 16439
rect 16807 16405 16816 16439
rect 16764 16396 16816 16405
rect 17316 16396 17368 16448
rect 21456 16464 21508 16516
rect 18144 16396 18196 16448
rect 18420 16396 18472 16448
rect 18512 16396 18564 16448
rect 19432 16396 19484 16448
rect 19616 16396 19668 16448
rect 20536 16439 20588 16448
rect 20536 16405 20545 16439
rect 20545 16405 20579 16439
rect 20579 16405 20588 16439
rect 20536 16396 20588 16405
rect 21824 16396 21876 16448
rect 24400 16464 24452 16516
rect 22652 16396 22704 16448
rect 3658 16294 3710 16346
rect 3722 16294 3774 16346
rect 3786 16294 3838 16346
rect 3850 16294 3902 16346
rect 3914 16294 3966 16346
rect 3978 16294 4030 16346
rect 7658 16294 7710 16346
rect 7722 16294 7774 16346
rect 7786 16294 7838 16346
rect 7850 16294 7902 16346
rect 7914 16294 7966 16346
rect 7978 16294 8030 16346
rect 11658 16294 11710 16346
rect 11722 16294 11774 16346
rect 11786 16294 11838 16346
rect 11850 16294 11902 16346
rect 11914 16294 11966 16346
rect 11978 16294 12030 16346
rect 15658 16294 15710 16346
rect 15722 16294 15774 16346
rect 15786 16294 15838 16346
rect 15850 16294 15902 16346
rect 15914 16294 15966 16346
rect 15978 16294 16030 16346
rect 19658 16294 19710 16346
rect 19722 16294 19774 16346
rect 19786 16294 19838 16346
rect 19850 16294 19902 16346
rect 19914 16294 19966 16346
rect 19978 16294 20030 16346
rect 23658 16294 23710 16346
rect 23722 16294 23774 16346
rect 23786 16294 23838 16346
rect 23850 16294 23902 16346
rect 23914 16294 23966 16346
rect 23978 16294 24030 16346
rect 2228 16124 2280 16176
rect 2136 16056 2188 16108
rect 4804 16192 4856 16244
rect 6644 16192 6696 16244
rect 7104 16192 7156 16244
rect 8208 16192 8260 16244
rect 4712 16124 4764 16176
rect 5172 16124 5224 16176
rect 5540 16124 5592 16176
rect 3792 16056 3844 16108
rect 5908 16099 5960 16108
rect 5908 16065 5917 16099
rect 5917 16065 5951 16099
rect 5951 16065 5960 16099
rect 5908 16056 5960 16065
rect 7288 16124 7340 16176
rect 8944 16124 8996 16176
rect 2780 15920 2832 15972
rect 5172 15988 5224 16040
rect 7564 16056 7616 16108
rect 4160 15920 4212 15972
rect 8300 16056 8352 16108
rect 10508 16192 10560 16244
rect 10692 16192 10744 16244
rect 10048 16124 10100 16176
rect 12624 16192 12676 16244
rect 14556 16192 14608 16244
rect 15568 16192 15620 16244
rect 16764 16192 16816 16244
rect 17316 16235 17368 16244
rect 17316 16201 17325 16235
rect 17325 16201 17359 16235
rect 17359 16201 17368 16235
rect 17316 16192 17368 16201
rect 17960 16192 18012 16244
rect 10324 16056 10376 16108
rect 9772 16031 9824 16040
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 10048 15988 10100 16040
rect 11428 16056 11480 16108
rect 3332 15852 3384 15904
rect 8116 15852 8168 15904
rect 9036 15895 9088 15904
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 10968 15988 11020 16040
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 11336 15963 11388 15972
rect 11336 15929 11345 15963
rect 11345 15929 11379 15963
rect 11379 15929 11388 15963
rect 11336 15920 11388 15929
rect 12624 15852 12676 15904
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 14280 16124 14332 16176
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 14004 15988 14056 16040
rect 15568 16056 15620 16108
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 16672 16099 16724 16108
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 16856 16099 16908 16108
rect 16856 16065 16863 16099
rect 16863 16065 16908 16099
rect 16856 16056 16908 16065
rect 14372 15988 14424 16040
rect 17224 16056 17276 16108
rect 18512 16235 18564 16244
rect 18512 16201 18521 16235
rect 18521 16201 18555 16235
rect 18555 16201 18564 16235
rect 18512 16192 18564 16201
rect 18972 16192 19024 16244
rect 19340 16192 19392 16244
rect 20352 16192 20404 16244
rect 22836 16192 22888 16244
rect 17408 15988 17460 16040
rect 17868 15988 17920 16040
rect 18420 15988 18472 16040
rect 18788 16124 18840 16176
rect 20536 16124 20588 16176
rect 21824 16167 21876 16176
rect 21824 16133 21833 16167
rect 21833 16133 21867 16167
rect 21867 16133 21876 16167
rect 21824 16124 21876 16133
rect 22560 16124 22612 16176
rect 18788 15988 18840 16040
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 19340 16099 19392 16108
rect 19340 16065 19349 16099
rect 19349 16065 19383 16099
rect 19383 16065 19392 16099
rect 19340 16056 19392 16065
rect 19524 16056 19576 16108
rect 20168 16056 20220 16108
rect 21548 16099 21600 16108
rect 21548 16065 21557 16099
rect 21557 16065 21591 16099
rect 21591 16065 21600 16099
rect 21548 16056 21600 16065
rect 26148 16056 26200 16108
rect 16120 15920 16172 15972
rect 16856 15920 16908 15972
rect 17132 15920 17184 15972
rect 20444 15920 20496 15972
rect 21824 15920 21876 15972
rect 14832 15852 14884 15904
rect 18144 15852 18196 15904
rect 25964 15852 26016 15904
rect 26240 15852 26292 15904
rect 2918 15750 2970 15802
rect 2982 15750 3034 15802
rect 3046 15750 3098 15802
rect 3110 15750 3162 15802
rect 3174 15750 3226 15802
rect 3238 15750 3290 15802
rect 6918 15750 6970 15802
rect 6982 15750 7034 15802
rect 7046 15750 7098 15802
rect 7110 15750 7162 15802
rect 7174 15750 7226 15802
rect 7238 15750 7290 15802
rect 10918 15750 10970 15802
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 11238 15750 11290 15802
rect 14918 15750 14970 15802
rect 14982 15750 15034 15802
rect 15046 15750 15098 15802
rect 15110 15750 15162 15802
rect 15174 15750 15226 15802
rect 15238 15750 15290 15802
rect 18918 15750 18970 15802
rect 18982 15750 19034 15802
rect 19046 15750 19098 15802
rect 19110 15750 19162 15802
rect 19174 15750 19226 15802
rect 19238 15750 19290 15802
rect 22918 15750 22970 15802
rect 22982 15750 23034 15802
rect 23046 15750 23098 15802
rect 23110 15750 23162 15802
rect 23174 15750 23226 15802
rect 23238 15750 23290 15802
rect 3792 15691 3844 15700
rect 3792 15657 3801 15691
rect 3801 15657 3835 15691
rect 3835 15657 3844 15691
rect 3792 15648 3844 15657
rect 4252 15648 4304 15700
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 7380 15648 7432 15700
rect 9588 15648 9640 15700
rect 10324 15691 10376 15700
rect 10324 15657 10333 15691
rect 10333 15657 10367 15691
rect 10367 15657 10376 15691
rect 10324 15648 10376 15657
rect 13544 15648 13596 15700
rect 14188 15648 14240 15700
rect 16120 15648 16172 15700
rect 16488 15648 16540 15700
rect 20076 15648 20128 15700
rect 19340 15623 19392 15632
rect 5080 15512 5132 15564
rect 5540 15555 5592 15564
rect 5540 15521 5549 15555
rect 5549 15521 5583 15555
rect 5583 15521 5592 15555
rect 5540 15512 5592 15521
rect 11704 15512 11756 15564
rect 15568 15512 15620 15564
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 3332 15444 3384 15496
rect 4712 15444 4764 15496
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 5172 15487 5224 15496
rect 5172 15453 5181 15487
rect 5181 15453 5215 15487
rect 5215 15453 5224 15487
rect 5172 15444 5224 15453
rect 8116 15487 8168 15496
rect 8116 15453 8134 15487
rect 8134 15453 8168 15487
rect 8116 15444 8168 15453
rect 8484 15444 8536 15496
rect 9680 15444 9732 15496
rect 5908 15376 5960 15428
rect 4436 15308 4488 15360
rect 7104 15376 7156 15428
rect 9036 15376 9088 15428
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 8116 15308 8168 15360
rect 10508 15444 10560 15496
rect 9864 15376 9916 15428
rect 10876 15487 10928 15496
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 11336 15444 11388 15496
rect 14832 15444 14884 15496
rect 19340 15589 19349 15623
rect 19349 15589 19383 15623
rect 19383 15589 19392 15623
rect 19340 15580 19392 15589
rect 21180 15580 21232 15632
rect 21548 15580 21600 15632
rect 24676 15512 24728 15564
rect 26148 15512 26200 15564
rect 18512 15444 18564 15496
rect 12256 15376 12308 15428
rect 15476 15376 15528 15428
rect 18052 15376 18104 15428
rect 12072 15308 12124 15360
rect 14740 15308 14792 15360
rect 17868 15308 17920 15360
rect 17960 15308 18012 15360
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 23480 15444 23532 15496
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 20076 15376 20128 15428
rect 24584 15376 24636 15428
rect 25964 15376 26016 15428
rect 22836 15308 22888 15360
rect 25044 15308 25096 15360
rect 26332 15351 26384 15360
rect 26332 15317 26341 15351
rect 26341 15317 26375 15351
rect 26375 15317 26384 15351
rect 26332 15308 26384 15317
rect 3658 15206 3710 15258
rect 3722 15206 3774 15258
rect 3786 15206 3838 15258
rect 3850 15206 3902 15258
rect 3914 15206 3966 15258
rect 3978 15206 4030 15258
rect 7658 15206 7710 15258
rect 7722 15206 7774 15258
rect 7786 15206 7838 15258
rect 7850 15206 7902 15258
rect 7914 15206 7966 15258
rect 7978 15206 8030 15258
rect 11658 15206 11710 15258
rect 11722 15206 11774 15258
rect 11786 15206 11838 15258
rect 11850 15206 11902 15258
rect 11914 15206 11966 15258
rect 11978 15206 12030 15258
rect 15658 15206 15710 15258
rect 15722 15206 15774 15258
rect 15786 15206 15838 15258
rect 15850 15206 15902 15258
rect 15914 15206 15966 15258
rect 15978 15206 16030 15258
rect 19658 15206 19710 15258
rect 19722 15206 19774 15258
rect 19786 15206 19838 15258
rect 19850 15206 19902 15258
rect 19914 15206 19966 15258
rect 19978 15206 20030 15258
rect 23658 15206 23710 15258
rect 23722 15206 23774 15258
rect 23786 15206 23838 15258
rect 23850 15206 23902 15258
rect 23914 15206 23966 15258
rect 23978 15206 24030 15258
rect 2136 15147 2188 15156
rect 2136 15113 2145 15147
rect 2145 15113 2179 15147
rect 2179 15113 2188 15147
rect 2136 15104 2188 15113
rect 4344 15104 4396 15156
rect 5908 15147 5960 15156
rect 5908 15113 5917 15147
rect 5917 15113 5951 15147
rect 5951 15113 5960 15147
rect 5908 15104 5960 15113
rect 6920 15104 6972 15156
rect 7104 15104 7156 15156
rect 8208 15104 8260 15156
rect 9864 15147 9916 15156
rect 9864 15113 9873 15147
rect 9873 15113 9907 15147
rect 9907 15113 9916 15147
rect 9864 15104 9916 15113
rect 3332 15036 3384 15088
rect 4160 15036 4212 15088
rect 2780 14968 2832 15020
rect 8944 15036 8996 15088
rect 10324 15104 10376 15156
rect 10876 15104 10928 15156
rect 11060 15104 11112 15156
rect 11428 15104 11480 15156
rect 16856 15104 16908 15156
rect 18420 15104 18472 15156
rect 2228 14900 2280 14952
rect 4804 14943 4856 14952
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 4896 14943 4948 14952
rect 4896 14909 4905 14943
rect 4905 14909 4939 14943
rect 4939 14909 4948 14943
rect 4896 14900 4948 14909
rect 4344 14807 4396 14816
rect 4344 14773 4353 14807
rect 4353 14773 4387 14807
rect 4387 14773 4396 14807
rect 4344 14764 4396 14773
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7012 14968 7064 15020
rect 7748 15011 7800 15020
rect 7748 14977 7757 15011
rect 7757 14977 7791 15011
rect 7791 14977 7800 15011
rect 7748 14968 7800 14977
rect 8208 15011 8260 15020
rect 8208 14977 8217 15011
rect 8217 14977 8251 15011
rect 8251 14977 8260 15011
rect 8208 14968 8260 14977
rect 8484 15011 8536 15020
rect 8484 14977 8500 15011
rect 8500 14977 8534 15011
rect 8534 14977 8536 15011
rect 8760 15011 8812 15020
rect 8484 14968 8536 14977
rect 8760 14977 8794 15011
rect 8794 14977 8812 15011
rect 8760 14968 8812 14977
rect 9036 14968 9088 15020
rect 7472 14943 7524 14952
rect 7472 14909 7481 14943
rect 7481 14909 7515 14943
rect 7515 14909 7524 14943
rect 7472 14900 7524 14909
rect 7564 14832 7616 14884
rect 8484 14832 8536 14884
rect 14004 15079 14056 15088
rect 14004 15045 14013 15079
rect 14013 15045 14047 15079
rect 14047 15045 14056 15079
rect 14004 15036 14056 15045
rect 17868 15036 17920 15088
rect 18604 15036 18656 15088
rect 10600 14968 10652 15020
rect 19340 15147 19392 15156
rect 19340 15113 19349 15147
rect 19349 15113 19383 15147
rect 19383 15113 19392 15147
rect 19340 15104 19392 15113
rect 19340 14968 19392 15020
rect 20076 15104 20128 15156
rect 22836 15036 22888 15088
rect 24124 14968 24176 15020
rect 24676 14968 24728 15020
rect 17684 14832 17736 14884
rect 21824 14943 21876 14952
rect 21824 14909 21833 14943
rect 21833 14909 21867 14943
rect 21867 14909 21876 14943
rect 21824 14900 21876 14909
rect 24216 14900 24268 14952
rect 25964 14943 26016 14952
rect 25964 14909 25973 14943
rect 25973 14909 26007 14943
rect 26007 14909 26016 14943
rect 25964 14900 26016 14909
rect 20444 14832 20496 14884
rect 9772 14764 9824 14816
rect 14832 14764 14884 14816
rect 24676 14764 24728 14816
rect 25136 14807 25188 14816
rect 25136 14773 25145 14807
rect 25145 14773 25179 14807
rect 25179 14773 25188 14807
rect 25136 14764 25188 14773
rect 26424 14764 26476 14816
rect 2918 14662 2970 14714
rect 2982 14662 3034 14714
rect 3046 14662 3098 14714
rect 3110 14662 3162 14714
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 6918 14662 6970 14714
rect 6982 14662 7034 14714
rect 7046 14662 7098 14714
rect 7110 14662 7162 14714
rect 7174 14662 7226 14714
rect 7238 14662 7290 14714
rect 10918 14662 10970 14714
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 11238 14662 11290 14714
rect 14918 14662 14970 14714
rect 14982 14662 15034 14714
rect 15046 14662 15098 14714
rect 15110 14662 15162 14714
rect 15174 14662 15226 14714
rect 15238 14662 15290 14714
rect 18918 14662 18970 14714
rect 18982 14662 19034 14714
rect 19046 14662 19098 14714
rect 19110 14662 19162 14714
rect 19174 14662 19226 14714
rect 19238 14662 19290 14714
rect 22918 14662 22970 14714
rect 22982 14662 23034 14714
rect 23046 14662 23098 14714
rect 23110 14662 23162 14714
rect 23174 14662 23226 14714
rect 23238 14662 23290 14714
rect 3332 14560 3384 14612
rect 6276 14560 6328 14612
rect 6828 14560 6880 14612
rect 8208 14560 8260 14612
rect 13728 14560 13780 14612
rect 18788 14560 18840 14612
rect 19340 14603 19392 14612
rect 19340 14569 19349 14603
rect 19349 14569 19383 14603
rect 19383 14569 19392 14603
rect 19340 14560 19392 14569
rect 19432 14560 19484 14612
rect 6736 14492 6788 14544
rect 7472 14492 7524 14544
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 12072 14492 12124 14544
rect 12716 14424 12768 14476
rect 13452 14424 13504 14476
rect 13728 14424 13780 14476
rect 4344 14356 4396 14408
rect 9864 14356 9916 14408
rect 9772 14288 9824 14340
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 15108 14288 15160 14340
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 18696 14492 18748 14544
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 16672 14356 16724 14408
rect 16948 14356 17000 14408
rect 17592 14356 17644 14408
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 18880 14399 18932 14408
rect 18880 14365 18888 14399
rect 18888 14365 18922 14399
rect 18922 14365 18932 14399
rect 18880 14356 18932 14365
rect 21180 14467 21232 14476
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 23572 14424 23624 14476
rect 24676 14467 24728 14476
rect 24676 14433 24685 14467
rect 24685 14433 24719 14467
rect 24719 14433 24728 14467
rect 24676 14424 24728 14433
rect 14832 14220 14884 14272
rect 15476 14220 15528 14272
rect 18604 14331 18656 14340
rect 18604 14297 18613 14331
rect 18613 14297 18647 14331
rect 18647 14297 18656 14331
rect 18604 14288 18656 14297
rect 18788 14220 18840 14272
rect 23480 14356 23532 14408
rect 24124 14356 24176 14408
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 26424 14399 26476 14408
rect 26424 14365 26433 14399
rect 26433 14365 26467 14399
rect 26467 14365 26476 14399
rect 26424 14356 26476 14365
rect 25136 14288 25188 14340
rect 22284 14220 22336 14272
rect 24860 14220 24912 14272
rect 3658 14118 3710 14170
rect 3722 14118 3774 14170
rect 3786 14118 3838 14170
rect 3850 14118 3902 14170
rect 3914 14118 3966 14170
rect 3978 14118 4030 14170
rect 7658 14118 7710 14170
rect 7722 14118 7774 14170
rect 7786 14118 7838 14170
rect 7850 14118 7902 14170
rect 7914 14118 7966 14170
rect 7978 14118 8030 14170
rect 11658 14118 11710 14170
rect 11722 14118 11774 14170
rect 11786 14118 11838 14170
rect 11850 14118 11902 14170
rect 11914 14118 11966 14170
rect 11978 14118 12030 14170
rect 15658 14118 15710 14170
rect 15722 14118 15774 14170
rect 15786 14118 15838 14170
rect 15850 14118 15902 14170
rect 15914 14118 15966 14170
rect 15978 14118 16030 14170
rect 19658 14118 19710 14170
rect 19722 14118 19774 14170
rect 19786 14118 19838 14170
rect 19850 14118 19902 14170
rect 19914 14118 19966 14170
rect 19978 14118 20030 14170
rect 23658 14118 23710 14170
rect 23722 14118 23774 14170
rect 23786 14118 23838 14170
rect 23850 14118 23902 14170
rect 23914 14118 23966 14170
rect 23978 14118 24030 14170
rect 7380 13948 7432 14000
rect 9772 13812 9824 13864
rect 10692 13923 10744 13932
rect 10692 13889 10701 13923
rect 10701 13889 10735 13923
rect 10735 13889 10744 13923
rect 10692 13880 10744 13889
rect 14188 14016 14240 14068
rect 15108 14016 15160 14068
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 18880 14016 18932 14068
rect 14280 13948 14332 14000
rect 18052 13948 18104 14000
rect 18696 13948 18748 14000
rect 22284 13991 22336 14000
rect 22284 13957 22293 13991
rect 22293 13957 22327 13991
rect 22327 13957 22336 13991
rect 22284 13948 22336 13957
rect 22836 13948 22888 14000
rect 24952 13948 25004 14000
rect 26332 13948 26384 14000
rect 11428 13880 11480 13932
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 10416 13787 10468 13796
rect 10416 13753 10425 13787
rect 10425 13753 10459 13787
rect 10459 13753 10468 13787
rect 10416 13744 10468 13753
rect 12072 13923 12124 13932
rect 12072 13889 12081 13923
rect 12081 13889 12115 13923
rect 12115 13889 12124 13923
rect 12072 13880 12124 13889
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 14464 13880 14516 13932
rect 15752 13880 15804 13932
rect 19432 13880 19484 13932
rect 20076 13880 20128 13932
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 12256 13812 12308 13864
rect 13544 13744 13596 13796
rect 4804 13676 4856 13728
rect 5264 13676 5316 13728
rect 11336 13676 11388 13728
rect 12532 13676 12584 13728
rect 13820 13676 13872 13728
rect 14372 13676 14424 13728
rect 16856 13744 16908 13796
rect 17316 13744 17368 13796
rect 18420 13744 18472 13796
rect 19340 13812 19392 13864
rect 20720 13812 20772 13864
rect 21824 13812 21876 13864
rect 22008 13855 22060 13864
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 22008 13812 22060 13821
rect 23480 13812 23532 13864
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 15844 13676 15896 13728
rect 16948 13676 17000 13728
rect 19524 13676 19576 13728
rect 25228 13676 25280 13728
rect 26148 13719 26200 13728
rect 26148 13685 26157 13719
rect 26157 13685 26191 13719
rect 26191 13685 26200 13719
rect 26148 13676 26200 13685
rect 2918 13574 2970 13626
rect 2982 13574 3034 13626
rect 3046 13574 3098 13626
rect 3110 13574 3162 13626
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 6918 13574 6970 13626
rect 6982 13574 7034 13626
rect 7046 13574 7098 13626
rect 7110 13574 7162 13626
rect 7174 13574 7226 13626
rect 7238 13574 7290 13626
rect 10918 13574 10970 13626
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 11238 13574 11290 13626
rect 14918 13574 14970 13626
rect 14982 13574 15034 13626
rect 15046 13574 15098 13626
rect 15110 13574 15162 13626
rect 15174 13574 15226 13626
rect 15238 13574 15290 13626
rect 18918 13574 18970 13626
rect 18982 13574 19034 13626
rect 19046 13574 19098 13626
rect 19110 13574 19162 13626
rect 19174 13574 19226 13626
rect 19238 13574 19290 13626
rect 22918 13574 22970 13626
rect 22982 13574 23034 13626
rect 23046 13574 23098 13626
rect 23110 13574 23162 13626
rect 23174 13574 23226 13626
rect 23238 13574 23290 13626
rect 4068 13336 4120 13388
rect 4896 13404 4948 13456
rect 4436 13379 4488 13388
rect 4436 13345 4445 13379
rect 4445 13345 4479 13379
rect 4479 13345 4488 13379
rect 4436 13336 4488 13345
rect 4988 13336 5040 13388
rect 7564 13472 7616 13524
rect 11520 13472 11572 13524
rect 11796 13472 11848 13524
rect 15384 13472 15436 13524
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 16212 13472 16264 13524
rect 18420 13472 18472 13524
rect 18788 13472 18840 13524
rect 22836 13472 22888 13524
rect 7380 13404 7432 13456
rect 8300 13404 8352 13456
rect 8944 13404 8996 13456
rect 9496 13404 9548 13456
rect 2044 13268 2096 13320
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4528 13268 4580 13320
rect 4804 13268 4856 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 5908 13311 5960 13320
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 6184 13311 6236 13320
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 6184 13268 6236 13277
rect 7104 13336 7156 13388
rect 9588 13336 9640 13388
rect 9956 13336 10008 13388
rect 10600 13336 10652 13388
rect 10692 13268 10744 13320
rect 18604 13404 18656 13456
rect 19248 13447 19300 13456
rect 19248 13413 19257 13447
rect 19257 13413 19291 13447
rect 19291 13413 19300 13447
rect 19248 13404 19300 13413
rect 13820 13336 13872 13388
rect 12532 13311 12584 13320
rect 12532 13277 12550 13311
rect 12550 13277 12584 13311
rect 12532 13268 12584 13277
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 18236 13336 18288 13388
rect 15844 13268 15896 13320
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 2136 13132 2188 13184
rect 2780 13175 2832 13184
rect 2780 13141 2789 13175
rect 2789 13141 2823 13175
rect 2823 13141 2832 13175
rect 2780 13132 2832 13141
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 4804 13132 4856 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 8760 13132 8812 13184
rect 9864 13200 9916 13252
rect 11336 13200 11388 13252
rect 10508 13132 10560 13184
rect 11060 13132 11112 13184
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 14188 13200 14240 13252
rect 16672 13268 16724 13320
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 18052 13268 18104 13320
rect 22008 13336 22060 13388
rect 25044 13379 25096 13388
rect 25044 13345 25053 13379
rect 25053 13345 25087 13379
rect 25087 13345 25096 13379
rect 25044 13336 25096 13345
rect 26240 13336 26292 13388
rect 20720 13268 20772 13320
rect 24124 13268 24176 13320
rect 18144 13200 18196 13252
rect 16764 13175 16816 13184
rect 16764 13141 16773 13175
rect 16773 13141 16807 13175
rect 16807 13141 16816 13175
rect 16764 13132 16816 13141
rect 18512 13132 18564 13184
rect 19340 13200 19392 13252
rect 25780 13132 25832 13184
rect 3658 13030 3710 13082
rect 3722 13030 3774 13082
rect 3786 13030 3838 13082
rect 3850 13030 3902 13082
rect 3914 13030 3966 13082
rect 3978 13030 4030 13082
rect 7658 13030 7710 13082
rect 7722 13030 7774 13082
rect 7786 13030 7838 13082
rect 7850 13030 7902 13082
rect 7914 13030 7966 13082
rect 7978 13030 8030 13082
rect 11658 13030 11710 13082
rect 11722 13030 11774 13082
rect 11786 13030 11838 13082
rect 11850 13030 11902 13082
rect 11914 13030 11966 13082
rect 11978 13030 12030 13082
rect 15658 13030 15710 13082
rect 15722 13030 15774 13082
rect 15786 13030 15838 13082
rect 15850 13030 15902 13082
rect 15914 13030 15966 13082
rect 15978 13030 16030 13082
rect 19658 13030 19710 13082
rect 19722 13030 19774 13082
rect 19786 13030 19838 13082
rect 19850 13030 19902 13082
rect 19914 13030 19966 13082
rect 19978 13030 20030 13082
rect 23658 13030 23710 13082
rect 23722 13030 23774 13082
rect 23786 13030 23838 13082
rect 23850 13030 23902 13082
rect 23914 13030 23966 13082
rect 23978 13030 24030 13082
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 2964 12928 3016 12980
rect 2780 12860 2832 12912
rect 848 12792 900 12844
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 4804 12928 4856 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 5540 12860 5592 12912
rect 6368 12860 6420 12912
rect 6736 12860 6788 12912
rect 6920 12860 6972 12912
rect 7380 12860 7432 12912
rect 5448 12792 5500 12844
rect 4068 12588 4120 12640
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 4712 12724 4764 12776
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 5448 12656 5500 12708
rect 7656 12792 7708 12844
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 10692 12928 10744 12980
rect 11520 12928 11572 12980
rect 12164 12928 12216 12980
rect 14464 12928 14516 12980
rect 15384 12928 15436 12980
rect 16488 12928 16540 12980
rect 9220 12860 9272 12912
rect 5632 12767 5684 12776
rect 5632 12733 5641 12767
rect 5641 12733 5675 12767
rect 5675 12733 5684 12767
rect 5632 12724 5684 12733
rect 6000 12724 6052 12776
rect 8576 12792 8628 12844
rect 9956 12792 10008 12844
rect 10232 12792 10284 12844
rect 11060 12835 11112 12844
rect 11060 12801 11078 12835
rect 11078 12801 11112 12835
rect 11060 12792 11112 12801
rect 8300 12724 8352 12776
rect 8484 12767 8536 12776
rect 8484 12733 8493 12767
rect 8493 12733 8527 12767
rect 8527 12733 8536 12767
rect 8484 12724 8536 12733
rect 4804 12588 4856 12640
rect 7564 12656 7616 12708
rect 11520 12724 11572 12776
rect 13084 12860 13136 12912
rect 14832 12903 14884 12912
rect 14832 12869 14841 12903
rect 14841 12869 14875 12903
rect 14875 12869 14884 12903
rect 14832 12860 14884 12869
rect 16764 12860 16816 12912
rect 18052 12971 18104 12980
rect 18052 12937 18061 12971
rect 18061 12937 18095 12971
rect 18095 12937 18104 12971
rect 18052 12928 18104 12937
rect 18512 12971 18564 12980
rect 18512 12937 18521 12971
rect 18521 12937 18555 12971
rect 18555 12937 18564 12971
rect 18512 12928 18564 12937
rect 18696 12928 18748 12980
rect 19248 12928 19300 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 20076 12928 20128 12980
rect 24400 12928 24452 12980
rect 19524 12860 19576 12912
rect 26148 12860 26200 12912
rect 9864 12631 9916 12640
rect 9864 12597 9873 12631
rect 9873 12597 9907 12631
rect 9907 12597 9916 12631
rect 9864 12588 9916 12597
rect 10232 12588 10284 12640
rect 14096 12792 14148 12844
rect 14924 12767 14976 12776
rect 14924 12733 14933 12767
rect 14933 12733 14967 12767
rect 14967 12733 14976 12767
rect 14924 12724 14976 12733
rect 14004 12631 14056 12640
rect 14004 12597 14013 12631
rect 14013 12597 14047 12631
rect 14047 12597 14056 12631
rect 14004 12588 14056 12597
rect 14832 12588 14884 12640
rect 18052 12724 18104 12776
rect 18236 12724 18288 12776
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 24952 12792 25004 12844
rect 17960 12656 18012 12708
rect 19432 12724 19484 12776
rect 18788 12588 18840 12640
rect 21180 12588 21232 12640
rect 24584 12631 24636 12640
rect 24584 12597 24593 12631
rect 24593 12597 24627 12631
rect 24627 12597 24636 12631
rect 24584 12588 24636 12597
rect 2918 12486 2970 12538
rect 2982 12486 3034 12538
rect 3046 12486 3098 12538
rect 3110 12486 3162 12538
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 6918 12486 6970 12538
rect 6982 12486 7034 12538
rect 7046 12486 7098 12538
rect 7110 12486 7162 12538
rect 7174 12486 7226 12538
rect 7238 12486 7290 12538
rect 10918 12486 10970 12538
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 11238 12486 11290 12538
rect 14918 12486 14970 12538
rect 14982 12486 15034 12538
rect 15046 12486 15098 12538
rect 15110 12486 15162 12538
rect 15174 12486 15226 12538
rect 15238 12486 15290 12538
rect 18918 12486 18970 12538
rect 18982 12486 19034 12538
rect 19046 12486 19098 12538
rect 19110 12486 19162 12538
rect 19174 12486 19226 12538
rect 19238 12486 19290 12538
rect 22918 12486 22970 12538
rect 22982 12486 23034 12538
rect 23046 12486 23098 12538
rect 23110 12486 23162 12538
rect 23174 12486 23226 12538
rect 23238 12486 23290 12538
rect 4160 12384 4212 12436
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 13268 12384 13320 12436
rect 19340 12384 19392 12436
rect 22192 12384 22244 12436
rect 10048 12316 10100 12368
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 8484 12248 8536 12300
rect 8944 12248 8996 12300
rect 10508 12248 10560 12300
rect 14740 12248 14792 12300
rect 20720 12248 20772 12300
rect 21180 12291 21232 12300
rect 21180 12257 21189 12291
rect 21189 12257 21223 12291
rect 21223 12257 21232 12291
rect 21180 12248 21232 12257
rect 24952 12291 25004 12300
rect 24952 12257 24961 12291
rect 24961 12257 24995 12291
rect 24995 12257 25004 12291
rect 24952 12248 25004 12257
rect 1584 12180 1636 12232
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 2136 12155 2188 12164
rect 2136 12121 2170 12155
rect 2170 12121 2188 12155
rect 2136 12112 2188 12121
rect 2320 12112 2372 12164
rect 5540 12180 5592 12232
rect 8760 12223 8812 12232
rect 8760 12189 8769 12223
rect 8769 12189 8803 12223
rect 8803 12189 8812 12223
rect 8760 12180 8812 12189
rect 18788 12223 18840 12232
rect 18788 12189 18797 12223
rect 18797 12189 18831 12223
rect 18831 12189 18840 12223
rect 18788 12180 18840 12189
rect 20812 12223 20864 12232
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 20812 12180 20864 12189
rect 22744 12180 22796 12232
rect 4620 12112 4672 12164
rect 6368 12112 6420 12164
rect 9404 12112 9456 12164
rect 4712 12044 4764 12096
rect 10692 12112 10744 12164
rect 14004 12112 14056 12164
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 12900 12044 12952 12096
rect 13360 12044 13412 12096
rect 20168 12044 20220 12096
rect 23572 12044 23624 12096
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 25780 12223 25832 12232
rect 25780 12189 25789 12223
rect 25789 12189 25823 12223
rect 25823 12189 25832 12223
rect 25780 12180 25832 12189
rect 24492 12044 24544 12096
rect 25780 12044 25832 12096
rect 3658 11942 3710 11994
rect 3722 11942 3774 11994
rect 3786 11942 3838 11994
rect 3850 11942 3902 11994
rect 3914 11942 3966 11994
rect 3978 11942 4030 11994
rect 7658 11942 7710 11994
rect 7722 11942 7774 11994
rect 7786 11942 7838 11994
rect 7850 11942 7902 11994
rect 7914 11942 7966 11994
rect 7978 11942 8030 11994
rect 11658 11942 11710 11994
rect 11722 11942 11774 11994
rect 11786 11942 11838 11994
rect 11850 11942 11902 11994
rect 11914 11942 11966 11994
rect 11978 11942 12030 11994
rect 15658 11942 15710 11994
rect 15722 11942 15774 11994
rect 15786 11942 15838 11994
rect 15850 11942 15902 11994
rect 15914 11942 15966 11994
rect 15978 11942 16030 11994
rect 19658 11942 19710 11994
rect 19722 11942 19774 11994
rect 19786 11942 19838 11994
rect 19850 11942 19902 11994
rect 19914 11942 19966 11994
rect 19978 11942 20030 11994
rect 23658 11942 23710 11994
rect 23722 11942 23774 11994
rect 23786 11942 23838 11994
rect 23850 11942 23902 11994
rect 23914 11942 23966 11994
rect 23978 11942 24030 11994
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 2136 11704 2188 11756
rect 4620 11883 4672 11892
rect 4620 11849 4629 11883
rect 4629 11849 4663 11883
rect 4663 11849 4672 11883
rect 4620 11840 4672 11849
rect 5908 11883 5960 11892
rect 5908 11849 5917 11883
rect 5917 11849 5951 11883
rect 5951 11849 5960 11883
rect 5908 11840 5960 11849
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 9680 11840 9732 11892
rect 9864 11840 9916 11892
rect 4528 11704 4580 11756
rect 4804 11747 4856 11756
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 6092 11704 6144 11756
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 10508 11772 10560 11824
rect 12256 11840 12308 11892
rect 20996 11840 21048 11892
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 22192 11840 22244 11892
rect 22744 11840 22796 11892
rect 10692 11815 10744 11824
rect 10692 11781 10701 11815
rect 10701 11781 10735 11815
rect 10735 11781 10744 11815
rect 10692 11772 10744 11781
rect 20168 11815 20220 11824
rect 20168 11781 20177 11815
rect 20177 11781 20211 11815
rect 20211 11781 20220 11815
rect 20168 11772 20220 11781
rect 21732 11772 21784 11824
rect 23572 11772 23624 11824
rect 10324 11704 10376 11756
rect 11336 11704 11388 11756
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 3332 11636 3384 11688
rect 3700 11679 3752 11688
rect 3700 11645 3709 11679
rect 3709 11645 3743 11679
rect 3743 11645 3752 11679
rect 3700 11636 3752 11645
rect 9404 11636 9456 11688
rect 16672 11704 16724 11756
rect 21456 11636 21508 11688
rect 22468 11679 22520 11688
rect 22468 11645 22477 11679
rect 22477 11645 22511 11679
rect 22511 11645 22520 11679
rect 22468 11636 22520 11645
rect 2596 11568 2648 11620
rect 21364 11568 21416 11620
rect 23388 11679 23440 11688
rect 23388 11645 23397 11679
rect 23397 11645 23431 11679
rect 23431 11645 23440 11679
rect 23388 11636 23440 11645
rect 24952 11636 25004 11688
rect 24768 11568 24820 11620
rect 6368 11500 6420 11552
rect 14464 11500 14516 11552
rect 25688 11500 25740 11552
rect 2918 11398 2970 11450
rect 2982 11398 3034 11450
rect 3046 11398 3098 11450
rect 3110 11398 3162 11450
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 6918 11398 6970 11450
rect 6982 11398 7034 11450
rect 7046 11398 7098 11450
rect 7110 11398 7162 11450
rect 7174 11398 7226 11450
rect 7238 11398 7290 11450
rect 10918 11398 10970 11450
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 11238 11398 11290 11450
rect 14918 11398 14970 11450
rect 14982 11398 15034 11450
rect 15046 11398 15098 11450
rect 15110 11398 15162 11450
rect 15174 11398 15226 11450
rect 15238 11398 15290 11450
rect 18918 11398 18970 11450
rect 18982 11398 19034 11450
rect 19046 11398 19098 11450
rect 19110 11398 19162 11450
rect 19174 11398 19226 11450
rect 19238 11398 19290 11450
rect 22918 11398 22970 11450
rect 22982 11398 23034 11450
rect 23046 11398 23098 11450
rect 23110 11398 23162 11450
rect 23174 11398 23226 11450
rect 23238 11398 23290 11450
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 2596 11092 2648 11144
rect 8208 11092 8260 11144
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 12716 11160 12768 11212
rect 16304 11228 16356 11280
rect 17776 11160 17828 11212
rect 4160 10956 4212 11008
rect 5172 10956 5224 11008
rect 12164 11024 12216 11076
rect 13176 11024 13228 11076
rect 14740 11024 14792 11076
rect 16304 11024 16356 11076
rect 8116 10956 8168 11008
rect 9588 10999 9640 11008
rect 9588 10965 9597 10999
rect 9597 10965 9631 10999
rect 9631 10965 9640 10999
rect 9588 10956 9640 10965
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 12072 10956 12124 10965
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 12900 10956 12952 11008
rect 15200 10999 15252 11008
rect 15200 10965 15209 10999
rect 15209 10965 15243 10999
rect 15243 10965 15252 10999
rect 15200 10956 15252 10965
rect 20812 11339 20864 11348
rect 20812 11305 20821 11339
rect 20821 11305 20855 11339
rect 20855 11305 20864 11339
rect 20812 11296 20864 11305
rect 21732 11339 21784 11348
rect 21732 11305 21741 11339
rect 21741 11305 21775 11339
rect 21775 11305 21784 11339
rect 21732 11296 21784 11305
rect 26056 11296 26108 11348
rect 19524 11228 19576 11280
rect 18696 11092 18748 11144
rect 21364 11203 21416 11212
rect 21364 11169 21373 11203
rect 21373 11169 21407 11203
rect 21407 11169 21416 11203
rect 21364 11160 21416 11169
rect 21456 11160 21508 11212
rect 23388 11160 23440 11212
rect 20996 11092 21048 11144
rect 22100 11092 22152 11144
rect 22744 11092 22796 11144
rect 20168 11024 20220 11076
rect 20444 11024 20496 11076
rect 21548 11024 21600 11076
rect 24124 11024 24176 11076
rect 24676 11067 24728 11076
rect 24676 11033 24685 11067
rect 24685 11033 24719 11067
rect 24719 11033 24728 11067
rect 24676 11024 24728 11033
rect 25688 11024 25740 11076
rect 18236 10956 18288 11008
rect 18420 10999 18472 11008
rect 18420 10965 18429 10999
rect 18429 10965 18463 10999
rect 18463 10965 18472 10999
rect 18420 10956 18472 10965
rect 18880 10999 18932 11008
rect 18880 10965 18889 10999
rect 18889 10965 18923 10999
rect 18923 10965 18932 10999
rect 18880 10956 18932 10965
rect 3658 10854 3710 10906
rect 3722 10854 3774 10906
rect 3786 10854 3838 10906
rect 3850 10854 3902 10906
rect 3914 10854 3966 10906
rect 3978 10854 4030 10906
rect 7658 10854 7710 10906
rect 7722 10854 7774 10906
rect 7786 10854 7838 10906
rect 7850 10854 7902 10906
rect 7914 10854 7966 10906
rect 7978 10854 8030 10906
rect 11658 10854 11710 10906
rect 11722 10854 11774 10906
rect 11786 10854 11838 10906
rect 11850 10854 11902 10906
rect 11914 10854 11966 10906
rect 11978 10854 12030 10906
rect 15658 10854 15710 10906
rect 15722 10854 15774 10906
rect 15786 10854 15838 10906
rect 15850 10854 15902 10906
rect 15914 10854 15966 10906
rect 15978 10854 16030 10906
rect 19658 10854 19710 10906
rect 19722 10854 19774 10906
rect 19786 10854 19838 10906
rect 19850 10854 19902 10906
rect 19914 10854 19966 10906
rect 19978 10854 20030 10906
rect 23658 10854 23710 10906
rect 23722 10854 23774 10906
rect 23786 10854 23838 10906
rect 23850 10854 23902 10906
rect 23914 10854 23966 10906
rect 23978 10854 24030 10906
rect 2780 10684 2832 10736
rect 3424 10684 3476 10736
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 4988 10752 5040 10804
rect 5080 10659 5132 10668
rect 5080 10625 5087 10659
rect 5087 10625 5132 10659
rect 5080 10616 5132 10625
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5356 10616 5408 10668
rect 6736 10616 6788 10668
rect 7564 10752 7616 10804
rect 7380 10684 7432 10736
rect 4804 10548 4856 10600
rect 7196 10616 7248 10668
rect 8944 10684 8996 10736
rect 10048 10795 10100 10804
rect 10048 10761 10057 10795
rect 10057 10761 10091 10795
rect 10091 10761 10100 10795
rect 10048 10752 10100 10761
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 11428 10752 11480 10804
rect 8116 10616 8168 10668
rect 9404 10616 9456 10668
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 10508 10616 10560 10668
rect 10232 10548 10284 10600
rect 7196 10480 7248 10532
rect 7472 10480 7524 10532
rect 9496 10480 9548 10532
rect 1492 10412 1544 10464
rect 5908 10412 5960 10464
rect 6092 10412 6144 10464
rect 8300 10412 8352 10464
rect 9312 10412 9364 10464
rect 9588 10412 9640 10464
rect 13176 10752 13228 10804
rect 13452 10752 13504 10804
rect 16304 10795 16356 10804
rect 16304 10761 16313 10795
rect 16313 10761 16347 10795
rect 16347 10761 16356 10795
rect 16304 10752 16356 10761
rect 16764 10752 16816 10804
rect 17316 10752 17368 10804
rect 18420 10752 18472 10804
rect 15200 10727 15252 10736
rect 15200 10693 15234 10727
rect 15234 10693 15252 10727
rect 15200 10684 15252 10693
rect 24492 10752 24544 10804
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 26056 10752 26108 10804
rect 20260 10684 20312 10736
rect 21916 10684 21968 10736
rect 13176 10616 13228 10668
rect 13728 10616 13780 10668
rect 12900 10548 12952 10600
rect 14004 10616 14056 10668
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 14832 10616 14884 10668
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 17684 10659 17736 10668
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 25044 10684 25096 10736
rect 14740 10548 14792 10600
rect 21456 10548 21508 10600
rect 24952 10616 25004 10668
rect 25136 10548 25188 10600
rect 25412 10591 25464 10600
rect 25412 10557 25421 10591
rect 25421 10557 25455 10591
rect 25455 10557 25464 10591
rect 25412 10548 25464 10557
rect 13728 10412 13780 10464
rect 14648 10455 14700 10464
rect 14648 10421 14657 10455
rect 14657 10421 14691 10455
rect 14691 10421 14700 10455
rect 14648 10412 14700 10421
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 17224 10455 17276 10464
rect 17224 10421 17233 10455
rect 17233 10421 17267 10455
rect 17267 10421 17276 10455
rect 17224 10412 17276 10421
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 21732 10412 21784 10464
rect 2918 10310 2970 10362
rect 2982 10310 3034 10362
rect 3046 10310 3098 10362
rect 3110 10310 3162 10362
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 6918 10310 6970 10362
rect 6982 10310 7034 10362
rect 7046 10310 7098 10362
rect 7110 10310 7162 10362
rect 7174 10310 7226 10362
rect 7238 10310 7290 10362
rect 10918 10310 10970 10362
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 11238 10310 11290 10362
rect 14918 10310 14970 10362
rect 14982 10310 15034 10362
rect 15046 10310 15098 10362
rect 15110 10310 15162 10362
rect 15174 10310 15226 10362
rect 15238 10310 15290 10362
rect 18918 10310 18970 10362
rect 18982 10310 19034 10362
rect 19046 10310 19098 10362
rect 19110 10310 19162 10362
rect 19174 10310 19226 10362
rect 19238 10310 19290 10362
rect 22918 10310 22970 10362
rect 22982 10310 23034 10362
rect 23046 10310 23098 10362
rect 23110 10310 23162 10362
rect 23174 10310 23226 10362
rect 23238 10310 23290 10362
rect 3332 10208 3384 10260
rect 4528 10208 4580 10260
rect 5356 10208 5408 10260
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 4160 10140 4212 10192
rect 4436 10140 4488 10192
rect 5448 10140 5500 10192
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 2780 10004 2832 10056
rect 3332 10004 3384 10056
rect 3792 10004 3844 10056
rect 5172 10072 5224 10124
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 7564 10208 7616 10260
rect 8208 10208 8260 10260
rect 6000 10140 6052 10192
rect 6736 10140 6788 10192
rect 1860 9868 1912 9920
rect 2780 9868 2832 9920
rect 3976 9868 4028 9920
rect 5080 10004 5132 10056
rect 5264 9936 5316 9988
rect 7104 10072 7156 10124
rect 7196 10115 7248 10124
rect 7196 10081 7205 10115
rect 7205 10081 7239 10115
rect 7239 10081 7248 10115
rect 7196 10072 7248 10081
rect 5816 9979 5868 9988
rect 5816 9945 5825 9979
rect 5825 9945 5859 9979
rect 5859 9945 5868 9979
rect 5816 9936 5868 9945
rect 5908 9936 5960 9988
rect 6368 10004 6420 10056
rect 7564 10004 7616 10056
rect 8300 10047 8352 10056
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 8576 10004 8628 10056
rect 10324 10208 10376 10260
rect 10416 10208 10468 10260
rect 12716 10208 12768 10260
rect 8944 10072 8996 10124
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 16396 10208 16448 10260
rect 16580 10208 16632 10260
rect 17408 10208 17460 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 17868 10208 17920 10260
rect 18880 10208 18932 10260
rect 25136 10251 25188 10260
rect 25136 10217 25145 10251
rect 25145 10217 25179 10251
rect 25179 10217 25188 10251
rect 25136 10208 25188 10217
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13820 10004 13872 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 4528 9911 4580 9920
rect 4528 9877 4537 9911
rect 4537 9877 4571 9911
rect 4571 9877 4580 9911
rect 4528 9868 4580 9877
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 5356 9868 5408 9920
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 5448 9868 5500 9877
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 7380 9936 7432 9988
rect 8116 9868 8168 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 8668 9868 8720 9920
rect 12072 9936 12124 9988
rect 13636 9936 13688 9988
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 14832 10115 14884 10124
rect 14832 10081 14841 10115
rect 14841 10081 14875 10115
rect 14875 10081 14884 10115
rect 14832 10072 14884 10081
rect 17684 10072 17736 10124
rect 21456 10115 21508 10124
rect 15292 9936 15344 9988
rect 16396 10004 16448 10056
rect 16672 10047 16724 10056
rect 16672 10013 16681 10047
rect 16681 10013 16715 10047
rect 16715 10013 16724 10047
rect 16672 10004 16724 10013
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 17040 10004 17092 10013
rect 16488 9979 16540 9988
rect 16488 9945 16497 9979
rect 16497 9945 16531 9979
rect 16531 9945 16540 9979
rect 16488 9936 16540 9945
rect 17408 10004 17460 10056
rect 18328 10004 18380 10056
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 21732 10115 21784 10124
rect 21732 10081 21741 10115
rect 21741 10081 21775 10115
rect 21775 10081 21784 10115
rect 21732 10072 21784 10081
rect 24124 10004 24176 10056
rect 24768 10004 24820 10056
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 25044 10047 25096 10056
rect 25044 10013 25053 10047
rect 25053 10013 25087 10047
rect 25087 10013 25096 10047
rect 25044 10004 25096 10013
rect 25228 10004 25280 10056
rect 25688 10004 25740 10056
rect 26148 10004 26200 10056
rect 12440 9868 12492 9920
rect 16212 9911 16264 9920
rect 16212 9877 16221 9911
rect 16221 9877 16255 9911
rect 16255 9877 16264 9911
rect 16212 9868 16264 9877
rect 18788 9979 18840 9988
rect 18788 9945 18806 9979
rect 18806 9945 18840 9979
rect 18788 9936 18840 9945
rect 18420 9868 18472 9920
rect 23296 9868 23348 9920
rect 24952 9911 25004 9920
rect 24952 9877 24961 9911
rect 24961 9877 24995 9911
rect 24995 9877 25004 9911
rect 24952 9868 25004 9877
rect 26332 9911 26384 9920
rect 26332 9877 26341 9911
rect 26341 9877 26375 9911
rect 26375 9877 26384 9911
rect 26332 9868 26384 9877
rect 3658 9766 3710 9818
rect 3722 9766 3774 9818
rect 3786 9766 3838 9818
rect 3850 9766 3902 9818
rect 3914 9766 3966 9818
rect 3978 9766 4030 9818
rect 7658 9766 7710 9818
rect 7722 9766 7774 9818
rect 7786 9766 7838 9818
rect 7850 9766 7902 9818
rect 7914 9766 7966 9818
rect 7978 9766 8030 9818
rect 11658 9766 11710 9818
rect 11722 9766 11774 9818
rect 11786 9766 11838 9818
rect 11850 9766 11902 9818
rect 11914 9766 11966 9818
rect 11978 9766 12030 9818
rect 15658 9766 15710 9818
rect 15722 9766 15774 9818
rect 15786 9766 15838 9818
rect 15850 9766 15902 9818
rect 15914 9766 15966 9818
rect 15978 9766 16030 9818
rect 19658 9766 19710 9818
rect 19722 9766 19774 9818
rect 19786 9766 19838 9818
rect 19850 9766 19902 9818
rect 19914 9766 19966 9818
rect 19978 9766 20030 9818
rect 23658 9766 23710 9818
rect 23722 9766 23774 9818
rect 23786 9766 23838 9818
rect 23850 9766 23902 9818
rect 23914 9766 23966 9818
rect 23978 9766 24030 9818
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 5264 9664 5316 9716
rect 5356 9664 5408 9716
rect 6828 9664 6880 9716
rect 7564 9664 7616 9716
rect 8116 9664 8168 9716
rect 10140 9664 10192 9716
rect 10416 9664 10468 9716
rect 14556 9664 14608 9716
rect 15292 9707 15344 9716
rect 15292 9673 15301 9707
rect 15301 9673 15335 9707
rect 15335 9673 15344 9707
rect 15292 9664 15344 9673
rect 16212 9664 16264 9716
rect 17040 9664 17092 9716
rect 18420 9707 18472 9716
rect 18420 9673 18429 9707
rect 18429 9673 18463 9707
rect 18463 9673 18472 9707
rect 18420 9664 18472 9673
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 5540 9596 5592 9648
rect 1492 9460 1544 9512
rect 2688 9528 2740 9580
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 4068 9528 4120 9580
rect 5172 9528 5224 9580
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 7472 9596 7524 9648
rect 12164 9596 12216 9648
rect 7380 9528 7432 9580
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 10600 9528 10652 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 14372 9571 14424 9580
rect 14372 9537 14381 9571
rect 14381 9537 14415 9571
rect 14415 9537 14424 9571
rect 14372 9528 14424 9537
rect 9220 9460 9272 9512
rect 10140 9460 10192 9512
rect 10324 9392 10376 9444
rect 10692 9392 10744 9444
rect 13452 9460 13504 9512
rect 11336 9392 11388 9444
rect 11428 9324 11480 9376
rect 16396 9528 16448 9580
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 18236 9596 18288 9648
rect 21916 9639 21968 9648
rect 21916 9605 21925 9639
rect 21925 9605 21959 9639
rect 21959 9605 21968 9639
rect 21916 9596 21968 9605
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 17592 9528 17644 9580
rect 17868 9528 17920 9580
rect 18052 9528 18104 9580
rect 18420 9528 18472 9580
rect 22836 9528 22888 9580
rect 24584 9528 24636 9580
rect 16856 9460 16908 9512
rect 19340 9460 19392 9512
rect 18696 9392 18748 9444
rect 17500 9324 17552 9376
rect 18052 9324 18104 9376
rect 22468 9460 22520 9512
rect 24216 9460 24268 9512
rect 26332 9596 26384 9648
rect 25228 9571 25280 9580
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 25688 9528 25740 9580
rect 25780 9571 25832 9580
rect 25780 9537 25789 9571
rect 25789 9537 25823 9571
rect 25823 9537 25832 9571
rect 25780 9528 25832 9537
rect 22100 9324 22152 9376
rect 22652 9324 22704 9376
rect 23940 9324 23992 9376
rect 25596 9324 25648 9376
rect 25780 9367 25832 9376
rect 25780 9333 25789 9367
rect 25789 9333 25823 9367
rect 25823 9333 25832 9367
rect 25780 9324 25832 9333
rect 2918 9222 2970 9274
rect 2982 9222 3034 9274
rect 3046 9222 3098 9274
rect 3110 9222 3162 9274
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 6918 9222 6970 9274
rect 6982 9222 7034 9274
rect 7046 9222 7098 9274
rect 7110 9222 7162 9274
rect 7174 9222 7226 9274
rect 7238 9222 7290 9274
rect 10918 9222 10970 9274
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 11238 9222 11290 9274
rect 14918 9222 14970 9274
rect 14982 9222 15034 9274
rect 15046 9222 15098 9274
rect 15110 9222 15162 9274
rect 15174 9222 15226 9274
rect 15238 9222 15290 9274
rect 18918 9222 18970 9274
rect 18982 9222 19034 9274
rect 19046 9222 19098 9274
rect 19110 9222 19162 9274
rect 19174 9222 19226 9274
rect 19238 9222 19290 9274
rect 22918 9222 22970 9274
rect 22982 9222 23034 9274
rect 23046 9222 23098 9274
rect 23110 9222 23162 9274
rect 23174 9222 23226 9274
rect 23238 9222 23290 9274
rect 2688 9120 2740 9172
rect 5080 9120 5132 9172
rect 7472 9120 7524 9172
rect 12440 9120 12492 9172
rect 3424 9052 3476 9104
rect 9680 9052 9732 9104
rect 14188 9120 14240 9172
rect 17408 9120 17460 9172
rect 18052 9120 18104 9172
rect 3516 8984 3568 9036
rect 9220 8984 9272 9036
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 1676 8848 1728 8900
rect 2780 8916 2832 8968
rect 4988 8916 5040 8968
rect 5540 8916 5592 8968
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 6368 8848 6420 8900
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 8760 8780 8812 8832
rect 10784 8780 10836 8832
rect 11428 8780 11480 8832
rect 12440 8780 12492 8832
rect 12624 8916 12676 8968
rect 16488 9052 16540 9104
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 12808 8848 12860 8900
rect 13268 8891 13320 8900
rect 13268 8857 13277 8891
rect 13277 8857 13311 8891
rect 13311 8857 13320 8891
rect 13268 8848 13320 8857
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 15384 8916 15436 8968
rect 17316 8916 17368 8968
rect 23572 9120 23624 9172
rect 24952 9120 25004 9172
rect 21456 9027 21508 9036
rect 21456 8993 21465 9027
rect 21465 8993 21499 9027
rect 21499 8993 21508 9027
rect 21456 8984 21508 8993
rect 23388 8984 23440 9036
rect 21640 8916 21692 8968
rect 22560 8916 22612 8968
rect 23664 8959 23716 8968
rect 23664 8925 23674 8959
rect 23674 8925 23708 8959
rect 23708 8925 23716 8959
rect 24860 8984 24912 9036
rect 25136 9095 25188 9104
rect 25136 9061 25145 9095
rect 25145 9061 25179 9095
rect 25179 9061 25188 9095
rect 25136 9052 25188 9061
rect 23664 8916 23716 8925
rect 23940 8959 23992 8968
rect 23940 8925 23949 8959
rect 23949 8925 23983 8959
rect 23983 8925 23992 8959
rect 23940 8916 23992 8925
rect 24124 8916 24176 8968
rect 16580 8848 16632 8900
rect 20720 8891 20772 8900
rect 20720 8857 20729 8891
rect 20729 8857 20763 8891
rect 20763 8857 20772 8891
rect 20720 8848 20772 8857
rect 21272 8848 21324 8900
rect 23480 8848 23532 8900
rect 24768 8916 24820 8968
rect 13820 8780 13872 8832
rect 14556 8780 14608 8832
rect 16488 8780 16540 8832
rect 17960 8780 18012 8832
rect 23572 8780 23624 8832
rect 24952 8848 25004 8900
rect 25780 8984 25832 9036
rect 25596 8959 25648 8968
rect 25596 8925 25605 8959
rect 25605 8925 25639 8959
rect 25639 8925 25648 8959
rect 25596 8916 25648 8925
rect 25780 8823 25832 8832
rect 25780 8789 25789 8823
rect 25789 8789 25823 8823
rect 25823 8789 25832 8823
rect 25780 8780 25832 8789
rect 3658 8678 3710 8730
rect 3722 8678 3774 8730
rect 3786 8678 3838 8730
rect 3850 8678 3902 8730
rect 3914 8678 3966 8730
rect 3978 8678 4030 8730
rect 7658 8678 7710 8730
rect 7722 8678 7774 8730
rect 7786 8678 7838 8730
rect 7850 8678 7902 8730
rect 7914 8678 7966 8730
rect 7978 8678 8030 8730
rect 11658 8678 11710 8730
rect 11722 8678 11774 8730
rect 11786 8678 11838 8730
rect 11850 8678 11902 8730
rect 11914 8678 11966 8730
rect 11978 8678 12030 8730
rect 15658 8678 15710 8730
rect 15722 8678 15774 8730
rect 15786 8678 15838 8730
rect 15850 8678 15902 8730
rect 15914 8678 15966 8730
rect 15978 8678 16030 8730
rect 19658 8678 19710 8730
rect 19722 8678 19774 8730
rect 19786 8678 19838 8730
rect 19850 8678 19902 8730
rect 19914 8678 19966 8730
rect 19978 8678 20030 8730
rect 23658 8678 23710 8730
rect 23722 8678 23774 8730
rect 23786 8678 23838 8730
rect 23850 8678 23902 8730
rect 23914 8678 23966 8730
rect 23978 8678 24030 8730
rect 5172 8551 5224 8560
rect 5172 8517 5181 8551
rect 5181 8517 5215 8551
rect 5215 8517 5224 8551
rect 5172 8508 5224 8517
rect 10508 8619 10560 8628
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 7380 8440 7432 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 8944 8440 8996 8492
rect 12808 8508 12860 8560
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 5908 8372 5960 8424
rect 6460 8372 6512 8424
rect 12164 8440 12216 8492
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 11428 8372 11480 8424
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 13820 8576 13872 8628
rect 14372 8576 14424 8628
rect 14556 8576 14608 8628
rect 14832 8508 14884 8560
rect 17408 8576 17460 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 13360 8483 13412 8492
rect 13360 8449 13394 8483
rect 13394 8449 13412 8483
rect 13360 8440 13412 8449
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 16396 8440 16448 8492
rect 20536 8576 20588 8628
rect 21548 8619 21600 8628
rect 21548 8585 21557 8619
rect 21557 8585 21591 8619
rect 21591 8585 21600 8619
rect 21548 8576 21600 8585
rect 24124 8576 24176 8628
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 21916 8508 21968 8560
rect 19800 8372 19852 8424
rect 19984 8372 20036 8424
rect 20168 8372 20220 8424
rect 21456 8440 21508 8492
rect 21640 8483 21692 8492
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 25136 8508 25188 8560
rect 22836 8440 22888 8492
rect 21088 8372 21140 8424
rect 21824 8372 21876 8424
rect 24124 8372 24176 8424
rect 7472 8236 7524 8288
rect 11704 8236 11756 8288
rect 13452 8236 13504 8288
rect 14556 8304 14608 8356
rect 15568 8347 15620 8356
rect 15568 8313 15577 8347
rect 15577 8313 15611 8347
rect 15611 8313 15620 8347
rect 15568 8304 15620 8313
rect 20536 8304 20588 8356
rect 20720 8304 20772 8356
rect 15476 8236 15528 8288
rect 15660 8236 15712 8288
rect 18604 8236 18656 8288
rect 21364 8236 21416 8288
rect 22192 8236 22244 8288
rect 22744 8279 22796 8288
rect 22744 8245 22753 8279
rect 22753 8245 22787 8279
rect 22787 8245 22796 8279
rect 22744 8236 22796 8245
rect 2918 8134 2970 8186
rect 2982 8134 3034 8186
rect 3046 8134 3098 8186
rect 3110 8134 3162 8186
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 6918 8134 6970 8186
rect 6982 8134 7034 8186
rect 7046 8134 7098 8186
rect 7110 8134 7162 8186
rect 7174 8134 7226 8186
rect 7238 8134 7290 8186
rect 10918 8134 10970 8186
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 11238 8134 11290 8186
rect 14918 8134 14970 8186
rect 14982 8134 15034 8186
rect 15046 8134 15098 8186
rect 15110 8134 15162 8186
rect 15174 8134 15226 8186
rect 15238 8134 15290 8186
rect 18918 8134 18970 8186
rect 18982 8134 19034 8186
rect 19046 8134 19098 8186
rect 19110 8134 19162 8186
rect 19174 8134 19226 8186
rect 19238 8134 19290 8186
rect 22918 8134 22970 8186
rect 22982 8134 23034 8186
rect 23046 8134 23098 8186
rect 23110 8134 23162 8186
rect 23174 8134 23226 8186
rect 23238 8134 23290 8186
rect 11428 8075 11480 8084
rect 11428 8041 11437 8075
rect 11437 8041 11471 8075
rect 11471 8041 11480 8075
rect 11428 8032 11480 8041
rect 12072 8032 12124 8084
rect 13360 8032 13412 8084
rect 14648 8032 14700 8084
rect 15660 8032 15712 8084
rect 15752 8032 15804 8084
rect 17132 8032 17184 8084
rect 17592 8075 17644 8084
rect 17592 8041 17601 8075
rect 17601 8041 17635 8075
rect 17635 8041 17644 8075
rect 17592 8032 17644 8041
rect 18236 8032 18288 8084
rect 20720 8032 20772 8084
rect 23572 8032 23624 8084
rect 13636 7964 13688 8016
rect 13728 7964 13780 8016
rect 8944 7896 8996 7948
rect 6460 7828 6512 7880
rect 7472 7828 7524 7880
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 11428 7896 11480 7948
rect 11612 7896 11664 7948
rect 4068 7760 4120 7812
rect 5540 7760 5592 7812
rect 8208 7760 8260 7812
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 11336 7828 11388 7880
rect 11704 7828 11756 7880
rect 13268 7828 13320 7880
rect 8116 7692 8168 7701
rect 10784 7735 10836 7744
rect 10784 7701 10793 7735
rect 10793 7701 10827 7735
rect 10827 7701 10836 7735
rect 14372 7828 14424 7880
rect 16120 7896 16172 7948
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 16488 7896 16540 7905
rect 16580 7896 16632 7948
rect 15476 7828 15528 7880
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 19708 7964 19760 8016
rect 20168 7964 20220 8016
rect 21824 7896 21876 7948
rect 21916 7939 21968 7948
rect 21916 7905 21925 7939
rect 21925 7905 21959 7939
rect 21959 7905 21968 7939
rect 21916 7896 21968 7905
rect 23296 7939 23348 7948
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 25964 7896 26016 7948
rect 14188 7760 14240 7812
rect 14556 7760 14608 7812
rect 14832 7760 14884 7812
rect 16580 7760 16632 7812
rect 19432 7828 19484 7880
rect 19800 7871 19852 7880
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 20076 7828 20128 7880
rect 20536 7828 20588 7880
rect 21180 7828 21232 7880
rect 21640 7828 21692 7880
rect 10784 7692 10836 7701
rect 15384 7692 15436 7744
rect 16212 7692 16264 7744
rect 19524 7760 19576 7812
rect 20444 7760 20496 7812
rect 20812 7760 20864 7812
rect 22192 7871 22244 7880
rect 22192 7837 22201 7871
rect 22201 7837 22235 7871
rect 22235 7837 22244 7871
rect 22192 7828 22244 7837
rect 22836 7828 22888 7880
rect 22468 7760 22520 7812
rect 24676 7760 24728 7812
rect 25780 7760 25832 7812
rect 3658 7590 3710 7642
rect 3722 7590 3774 7642
rect 3786 7590 3838 7642
rect 3850 7590 3902 7642
rect 3914 7590 3966 7642
rect 3978 7590 4030 7642
rect 7658 7590 7710 7642
rect 7722 7590 7774 7642
rect 7786 7590 7838 7642
rect 7850 7590 7902 7642
rect 7914 7590 7966 7642
rect 7978 7590 8030 7642
rect 11658 7590 11710 7642
rect 11722 7590 11774 7642
rect 11786 7590 11838 7642
rect 11850 7590 11902 7642
rect 11914 7590 11966 7642
rect 11978 7590 12030 7642
rect 15658 7590 15710 7642
rect 15722 7590 15774 7642
rect 15786 7590 15838 7642
rect 15850 7590 15902 7642
rect 15914 7590 15966 7642
rect 15978 7590 16030 7642
rect 19658 7590 19710 7642
rect 19722 7590 19774 7642
rect 19786 7590 19838 7642
rect 19850 7590 19902 7642
rect 19914 7590 19966 7642
rect 19978 7590 20030 7642
rect 23658 7590 23710 7642
rect 23722 7590 23774 7642
rect 23786 7590 23838 7642
rect 23850 7590 23902 7642
rect 23914 7590 23966 7642
rect 23978 7590 24030 7642
rect 2780 7488 2832 7540
rect 3516 7420 3568 7472
rect 4068 7463 4120 7472
rect 4068 7429 4077 7463
rect 4077 7429 4111 7463
rect 4111 7429 4120 7463
rect 4068 7420 4120 7429
rect 4528 7488 4580 7540
rect 5724 7488 5776 7540
rect 7380 7488 7432 7540
rect 8116 7488 8168 7540
rect 9128 7488 9180 7540
rect 10784 7488 10836 7540
rect 12624 7488 12676 7540
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 10140 7463 10192 7472
rect 10140 7429 10149 7463
rect 10149 7429 10183 7463
rect 10183 7429 10192 7463
rect 10140 7420 10192 7429
rect 12072 7463 12124 7472
rect 12072 7429 12106 7463
rect 12106 7429 12124 7463
rect 12072 7420 12124 7429
rect 14556 7488 14608 7540
rect 16764 7488 16816 7540
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 17592 7488 17644 7540
rect 19432 7488 19484 7540
rect 18420 7420 18472 7472
rect 18512 7420 18564 7472
rect 5448 7352 5500 7404
rect 7564 7352 7616 7404
rect 1860 7216 1912 7268
rect 3608 7284 3660 7336
rect 4620 7284 4672 7336
rect 6184 7284 6236 7336
rect 6828 7284 6880 7336
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 8024 7284 8076 7336
rect 8208 7395 8260 7404
rect 8208 7361 8218 7395
rect 8218 7361 8252 7395
rect 8252 7361 8260 7395
rect 8208 7352 8260 7361
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 8576 7395 8628 7404
rect 8576 7361 8590 7395
rect 8590 7361 8624 7395
rect 8624 7361 8628 7395
rect 8576 7352 8628 7361
rect 10600 7352 10652 7404
rect 10968 7352 11020 7404
rect 14004 7352 14056 7404
rect 10324 7327 10376 7336
rect 10324 7293 10333 7327
rect 10333 7293 10367 7327
rect 10367 7293 10376 7327
rect 10324 7284 10376 7293
rect 11520 7284 11572 7336
rect 13452 7284 13504 7336
rect 8300 7216 8352 7268
rect 11244 7216 11296 7268
rect 1676 7148 1728 7200
rect 5264 7148 5316 7200
rect 6736 7148 6788 7200
rect 8760 7191 8812 7200
rect 8760 7157 8769 7191
rect 8769 7157 8803 7191
rect 8803 7157 8812 7191
rect 8760 7148 8812 7157
rect 9956 7148 10008 7200
rect 10324 7148 10376 7200
rect 14096 7148 14148 7200
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 18604 7352 18656 7404
rect 17316 7327 17368 7336
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 17776 7284 17828 7336
rect 18696 7284 18748 7336
rect 19524 7352 19576 7404
rect 20076 7352 20128 7404
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 21272 7420 21324 7472
rect 25136 7488 25188 7540
rect 25412 7488 25464 7540
rect 26516 7531 26568 7540
rect 26516 7497 26525 7531
rect 26525 7497 26559 7531
rect 26559 7497 26568 7531
rect 26516 7488 26568 7497
rect 19708 7284 19760 7336
rect 20168 7284 20220 7336
rect 20720 7284 20772 7336
rect 21088 7284 21140 7336
rect 22376 7352 22428 7404
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 16396 7216 16448 7268
rect 21732 7284 21784 7336
rect 23572 7352 23624 7404
rect 24860 7352 24912 7404
rect 26332 7395 26384 7404
rect 26332 7361 26341 7395
rect 26341 7361 26375 7395
rect 26375 7361 26384 7395
rect 26332 7352 26384 7361
rect 18788 7148 18840 7200
rect 20352 7148 20404 7200
rect 20444 7148 20496 7200
rect 20904 7148 20956 7200
rect 21640 7259 21692 7268
rect 21640 7225 21649 7259
rect 21649 7225 21683 7259
rect 21683 7225 21692 7259
rect 21640 7216 21692 7225
rect 22376 7216 22428 7268
rect 22744 7216 22796 7268
rect 22100 7148 22152 7200
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 2918 7046 2970 7098
rect 2982 7046 3034 7098
rect 3046 7046 3098 7098
rect 3110 7046 3162 7098
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 6918 7046 6970 7098
rect 6982 7046 7034 7098
rect 7046 7046 7098 7098
rect 7110 7046 7162 7098
rect 7174 7046 7226 7098
rect 7238 7046 7290 7098
rect 10918 7046 10970 7098
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 11238 7046 11290 7098
rect 14918 7046 14970 7098
rect 14982 7046 15034 7098
rect 15046 7046 15098 7098
rect 15110 7046 15162 7098
rect 15174 7046 15226 7098
rect 15238 7046 15290 7098
rect 18918 7046 18970 7098
rect 18982 7046 19034 7098
rect 19046 7046 19098 7098
rect 19110 7046 19162 7098
rect 19174 7046 19226 7098
rect 19238 7046 19290 7098
rect 22918 7046 22970 7098
rect 22982 7046 23034 7098
rect 23046 7046 23098 7098
rect 23110 7046 23162 7098
rect 23174 7046 23226 7098
rect 23238 7046 23290 7098
rect 5172 6944 5224 6996
rect 6828 6944 6880 6996
rect 7564 6944 7616 6996
rect 8024 6944 8076 6996
rect 10784 6944 10836 6996
rect 11428 6944 11480 6996
rect 14648 6944 14700 6996
rect 8208 6876 8260 6928
rect 8300 6876 8352 6928
rect 8392 6876 8444 6928
rect 15384 6944 15436 6996
rect 16488 6944 16540 6996
rect 18788 6944 18840 6996
rect 19524 6944 19576 6996
rect 20444 6944 20496 6996
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 1860 6740 1912 6792
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 20904 6876 20956 6928
rect 21272 6876 21324 6928
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 5356 6783 5408 6792
rect 5356 6749 5366 6783
rect 5366 6749 5400 6783
rect 5400 6749 5408 6783
rect 5356 6740 5408 6749
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 3332 6647 3384 6656
rect 3332 6613 3341 6647
rect 3341 6613 3375 6647
rect 3375 6613 3384 6647
rect 3332 6604 3384 6613
rect 4712 6604 4764 6656
rect 6368 6740 6420 6792
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6736 6783 6788 6792
rect 6736 6749 6770 6783
rect 6770 6749 6788 6783
rect 6736 6740 6788 6749
rect 8208 6740 8260 6792
rect 8668 6740 8720 6792
rect 9864 6740 9916 6792
rect 14832 6740 14884 6792
rect 15568 6740 15620 6792
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 13544 6672 13596 6724
rect 16580 6672 16632 6724
rect 8116 6604 8168 6656
rect 9680 6604 9732 6656
rect 9772 6604 9824 6656
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 19708 6740 19760 6792
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 20720 6808 20772 6860
rect 21916 6944 21968 6996
rect 25228 6987 25280 6996
rect 25228 6953 25237 6987
rect 25237 6953 25271 6987
rect 25271 6953 25280 6987
rect 25228 6944 25280 6953
rect 19248 6672 19300 6724
rect 19432 6672 19484 6724
rect 20536 6740 20588 6792
rect 20628 6783 20680 6792
rect 20628 6749 20637 6783
rect 20637 6749 20671 6783
rect 20671 6749 20680 6783
rect 20628 6740 20680 6749
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 22100 6783 22152 6792
rect 22100 6749 22109 6783
rect 22109 6749 22143 6783
rect 22143 6749 22152 6783
rect 22100 6740 22152 6749
rect 22560 6740 22612 6792
rect 23112 6740 23164 6792
rect 23572 6740 23624 6792
rect 24216 6740 24268 6792
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 24952 6851 25004 6860
rect 24952 6817 24961 6851
rect 24961 6817 24995 6851
rect 24995 6817 25004 6851
rect 24952 6808 25004 6817
rect 25688 6851 25740 6860
rect 25688 6817 25697 6851
rect 25697 6817 25731 6851
rect 25731 6817 25740 6851
rect 25688 6808 25740 6817
rect 19340 6604 19392 6656
rect 20996 6647 21048 6656
rect 20996 6613 21005 6647
rect 21005 6613 21039 6647
rect 21039 6613 21048 6647
rect 20996 6604 21048 6613
rect 21548 6672 21600 6724
rect 22836 6715 22888 6724
rect 22836 6681 22845 6715
rect 22845 6681 22879 6715
rect 22879 6681 22888 6715
rect 22836 6672 22888 6681
rect 22192 6604 22244 6656
rect 22560 6604 22612 6656
rect 25320 6740 25372 6792
rect 25688 6672 25740 6724
rect 25504 6604 25556 6656
rect 25596 6604 25648 6656
rect 3658 6502 3710 6554
rect 3722 6502 3774 6554
rect 3786 6502 3838 6554
rect 3850 6502 3902 6554
rect 3914 6502 3966 6554
rect 3978 6502 4030 6554
rect 7658 6502 7710 6554
rect 7722 6502 7774 6554
rect 7786 6502 7838 6554
rect 7850 6502 7902 6554
rect 7914 6502 7966 6554
rect 7978 6502 8030 6554
rect 11658 6502 11710 6554
rect 11722 6502 11774 6554
rect 11786 6502 11838 6554
rect 11850 6502 11902 6554
rect 11914 6502 11966 6554
rect 11978 6502 12030 6554
rect 15658 6502 15710 6554
rect 15722 6502 15774 6554
rect 15786 6502 15838 6554
rect 15850 6502 15902 6554
rect 15914 6502 15966 6554
rect 15978 6502 16030 6554
rect 19658 6502 19710 6554
rect 19722 6502 19774 6554
rect 19786 6502 19838 6554
rect 19850 6502 19902 6554
rect 19914 6502 19966 6554
rect 19978 6502 20030 6554
rect 23658 6502 23710 6554
rect 23722 6502 23774 6554
rect 23786 6502 23838 6554
rect 23850 6502 23902 6554
rect 23914 6502 23966 6554
rect 23978 6502 24030 6554
rect 3424 6400 3476 6452
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 5448 6400 5500 6452
rect 8484 6400 8536 6452
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10232 6400 10284 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 13728 6400 13780 6452
rect 16212 6400 16264 6452
rect 18788 6400 18840 6452
rect 20168 6400 20220 6452
rect 20260 6400 20312 6452
rect 21640 6400 21692 6452
rect 21732 6400 21784 6452
rect 1860 6332 1912 6384
rect 3332 6332 3384 6384
rect 5356 6332 5408 6384
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 4528 6264 4580 6316
rect 6460 6332 6512 6384
rect 6828 6332 6880 6384
rect 8668 6332 8720 6384
rect 8760 6332 8812 6384
rect 6644 6307 6696 6316
rect 6644 6273 6678 6307
rect 6678 6273 6696 6307
rect 6644 6264 6696 6273
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 9496 6264 9548 6273
rect 9772 6307 9824 6316
rect 9772 6273 9806 6307
rect 9806 6273 9824 6307
rect 9772 6264 9824 6273
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 1400 6128 1452 6180
rect 1768 6060 1820 6112
rect 3516 6060 3568 6112
rect 7380 6196 7432 6248
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 17776 6332 17828 6384
rect 11796 6307 11848 6316
rect 11796 6273 11830 6307
rect 11830 6273 11848 6307
rect 11796 6264 11848 6273
rect 18604 6264 18656 6316
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 20536 6332 20588 6384
rect 20628 6332 20680 6384
rect 19432 6264 19484 6316
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 13544 6196 13596 6248
rect 16396 6196 16448 6248
rect 7564 6060 7616 6112
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 8852 6060 8904 6112
rect 12992 6103 13044 6112
rect 12992 6069 13001 6103
rect 13001 6069 13035 6103
rect 13035 6069 13044 6103
rect 12992 6060 13044 6069
rect 18788 6128 18840 6180
rect 19248 6128 19300 6180
rect 20720 6307 20772 6316
rect 20720 6273 20729 6307
rect 20729 6273 20763 6307
rect 20763 6273 20772 6307
rect 20720 6264 20772 6273
rect 20444 6196 20496 6248
rect 21548 6375 21600 6384
rect 21548 6341 21557 6375
rect 21557 6341 21591 6375
rect 21591 6341 21600 6375
rect 21548 6332 21600 6341
rect 23388 6400 23440 6452
rect 23572 6443 23624 6452
rect 23572 6409 23581 6443
rect 23581 6409 23615 6443
rect 23615 6409 23624 6443
rect 23572 6400 23624 6409
rect 21916 6264 21968 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 24860 6400 24912 6452
rect 25412 6443 25464 6452
rect 25412 6409 25437 6443
rect 25437 6409 25464 6443
rect 25412 6400 25464 6409
rect 22836 6307 22888 6316
rect 22836 6273 22845 6307
rect 22845 6273 22879 6307
rect 22879 6273 22888 6307
rect 22836 6264 22888 6273
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 22652 6196 22704 6248
rect 20904 6128 20956 6180
rect 19156 6060 19208 6112
rect 19432 6060 19484 6112
rect 19616 6060 19668 6112
rect 20812 6060 20864 6112
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 21916 6060 21968 6112
rect 22100 6060 22152 6112
rect 24032 6264 24084 6316
rect 24308 6332 24360 6384
rect 25228 6375 25280 6384
rect 24584 6264 24636 6316
rect 23940 6239 23992 6248
rect 23940 6205 23949 6239
rect 23949 6205 23983 6239
rect 23983 6205 23992 6239
rect 23940 6196 23992 6205
rect 25228 6341 25237 6375
rect 25237 6341 25271 6375
rect 25271 6341 25280 6375
rect 25228 6332 25280 6341
rect 24768 6307 24820 6316
rect 24768 6273 24777 6307
rect 24777 6273 24811 6307
rect 24811 6273 24820 6307
rect 24768 6264 24820 6273
rect 24860 6239 24912 6248
rect 24860 6205 24869 6239
rect 24869 6205 24903 6239
rect 24903 6205 24912 6239
rect 24860 6196 24912 6205
rect 24768 6128 24820 6180
rect 25596 6332 25648 6384
rect 25688 6307 25740 6316
rect 25688 6273 25697 6307
rect 25697 6273 25731 6307
rect 25731 6273 25740 6307
rect 25688 6264 25740 6273
rect 25964 6307 26016 6316
rect 25964 6273 25973 6307
rect 25973 6273 26007 6307
rect 26007 6273 26016 6307
rect 25964 6264 26016 6273
rect 24860 6060 24912 6112
rect 25320 6060 25372 6112
rect 25504 6128 25556 6180
rect 25596 6103 25648 6112
rect 25596 6069 25605 6103
rect 25605 6069 25639 6103
rect 25639 6069 25648 6103
rect 25596 6060 25648 6069
rect 26056 6103 26108 6112
rect 26056 6069 26065 6103
rect 26065 6069 26099 6103
rect 26099 6069 26108 6103
rect 26056 6060 26108 6069
rect 2918 5958 2970 6010
rect 2982 5958 3034 6010
rect 3046 5958 3098 6010
rect 3110 5958 3162 6010
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 6918 5958 6970 6010
rect 6982 5958 7034 6010
rect 7046 5958 7098 6010
rect 7110 5958 7162 6010
rect 7174 5958 7226 6010
rect 7238 5958 7290 6010
rect 10918 5958 10970 6010
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 11238 5958 11290 6010
rect 14918 5958 14970 6010
rect 14982 5958 15034 6010
rect 15046 5958 15098 6010
rect 15110 5958 15162 6010
rect 15174 5958 15226 6010
rect 15238 5958 15290 6010
rect 18918 5958 18970 6010
rect 18982 5958 19034 6010
rect 19046 5958 19098 6010
rect 19110 5958 19162 6010
rect 19174 5958 19226 6010
rect 19238 5958 19290 6010
rect 22918 5958 22970 6010
rect 22982 5958 23034 6010
rect 23046 5958 23098 6010
rect 23110 5958 23162 6010
rect 23174 5958 23226 6010
rect 23238 5958 23290 6010
rect 1952 5856 2004 5908
rect 2780 5856 2832 5908
rect 6644 5856 6696 5908
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 8668 5856 8720 5908
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 11796 5856 11848 5908
rect 4068 5788 4120 5840
rect 13176 5856 13228 5908
rect 16212 5856 16264 5908
rect 19432 5856 19484 5908
rect 23572 5856 23624 5908
rect 24768 5856 24820 5908
rect 12716 5788 12768 5840
rect 10692 5720 10744 5772
rect 16856 5788 16908 5840
rect 1768 5652 1820 5704
rect 7840 5652 7892 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 12992 5652 13044 5704
rect 13728 5652 13780 5704
rect 14004 5652 14056 5704
rect 16212 5763 16264 5772
rect 16212 5729 16221 5763
rect 16221 5729 16255 5763
rect 16255 5729 16264 5763
rect 16212 5720 16264 5729
rect 17132 5720 17184 5772
rect 18052 5652 18104 5704
rect 18696 5788 18748 5840
rect 19524 5720 19576 5772
rect 7564 5584 7616 5636
rect 13544 5584 13596 5636
rect 16672 5584 16724 5636
rect 18788 5652 18840 5704
rect 19616 5652 19668 5704
rect 20352 5788 20404 5840
rect 21180 5788 21232 5840
rect 20812 5720 20864 5772
rect 21732 5720 21784 5772
rect 22284 5720 22336 5772
rect 6368 5516 6420 5568
rect 8116 5516 8168 5568
rect 9404 5516 9456 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 16856 5516 16908 5568
rect 18604 5584 18656 5636
rect 18972 5584 19024 5636
rect 20076 5652 20128 5704
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 20996 5652 21048 5704
rect 21088 5695 21140 5704
rect 21088 5661 21097 5695
rect 21097 5661 21131 5695
rect 21131 5661 21140 5695
rect 21088 5652 21140 5661
rect 21180 5652 21232 5704
rect 20444 5584 20496 5636
rect 21824 5652 21876 5704
rect 22192 5652 22244 5704
rect 22560 5695 22612 5704
rect 22560 5661 22569 5695
rect 22569 5661 22603 5695
rect 22603 5661 22612 5695
rect 22560 5652 22612 5661
rect 25596 5788 25648 5840
rect 24860 5763 24912 5772
rect 24860 5729 24869 5763
rect 24869 5729 24903 5763
rect 24903 5729 24912 5763
rect 24860 5720 24912 5729
rect 25136 5720 25188 5772
rect 26056 5788 26108 5840
rect 24308 5652 24360 5704
rect 24768 5695 24820 5704
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 25228 5652 25280 5704
rect 25596 5695 25648 5704
rect 25596 5661 25605 5695
rect 25605 5661 25639 5695
rect 25639 5661 25648 5695
rect 25596 5652 25648 5661
rect 22192 5559 22244 5568
rect 22192 5525 22201 5559
rect 22201 5525 22235 5559
rect 22235 5525 22244 5559
rect 22192 5516 22244 5525
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 25228 5559 25280 5568
rect 25228 5525 25237 5559
rect 25237 5525 25271 5559
rect 25271 5525 25280 5559
rect 25228 5516 25280 5525
rect 3658 5414 3710 5466
rect 3722 5414 3774 5466
rect 3786 5414 3838 5466
rect 3850 5414 3902 5466
rect 3914 5414 3966 5466
rect 3978 5414 4030 5466
rect 7658 5414 7710 5466
rect 7722 5414 7774 5466
rect 7786 5414 7838 5466
rect 7850 5414 7902 5466
rect 7914 5414 7966 5466
rect 7978 5414 8030 5466
rect 11658 5414 11710 5466
rect 11722 5414 11774 5466
rect 11786 5414 11838 5466
rect 11850 5414 11902 5466
rect 11914 5414 11966 5466
rect 11978 5414 12030 5466
rect 15658 5414 15710 5466
rect 15722 5414 15774 5466
rect 15786 5414 15838 5466
rect 15850 5414 15902 5466
rect 15914 5414 15966 5466
rect 15978 5414 16030 5466
rect 19658 5414 19710 5466
rect 19722 5414 19774 5466
rect 19786 5414 19838 5466
rect 19850 5414 19902 5466
rect 19914 5414 19966 5466
rect 19978 5414 20030 5466
rect 23658 5414 23710 5466
rect 23722 5414 23774 5466
rect 23786 5414 23838 5466
rect 23850 5414 23902 5466
rect 23914 5414 23966 5466
rect 23978 5414 24030 5466
rect 8208 5312 8260 5364
rect 9036 5312 9088 5364
rect 7932 5287 7984 5296
rect 7932 5253 7941 5287
rect 7941 5253 7975 5287
rect 7975 5253 7984 5287
rect 7932 5244 7984 5253
rect 13268 5244 13320 5296
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 6000 5176 6052 5228
rect 4620 5151 4672 5160
rect 4620 5117 4629 5151
rect 4629 5117 4663 5151
rect 4663 5117 4672 5151
rect 4620 5108 4672 5117
rect 5172 5108 5224 5160
rect 8116 5219 8168 5228
rect 8116 5185 8130 5219
rect 8130 5185 8164 5219
rect 8164 5185 8168 5219
rect 8116 5176 8168 5185
rect 9772 5176 9824 5228
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 14096 5312 14148 5364
rect 14464 5312 14516 5364
rect 16396 5312 16448 5364
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 8300 5108 8352 5160
rect 9404 5108 9456 5160
rect 8208 5040 8260 5092
rect 13084 5108 13136 5160
rect 18420 5312 18472 5364
rect 19340 5244 19392 5296
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 17316 5176 17368 5228
rect 18696 5176 18748 5228
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 21088 5244 21140 5296
rect 20352 5176 20404 5228
rect 20444 5219 20496 5228
rect 20444 5185 20453 5219
rect 20453 5185 20487 5219
rect 20487 5185 20496 5219
rect 20444 5176 20496 5185
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 20812 5176 20864 5228
rect 14832 5108 14884 5160
rect 3976 4972 4028 5024
rect 4712 4972 4764 5024
rect 7472 4972 7524 5024
rect 18788 5040 18840 5092
rect 19984 5108 20036 5160
rect 20996 5108 21048 5160
rect 8944 4972 8996 5024
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 20168 5040 20220 5092
rect 20812 5040 20864 5092
rect 2918 4870 2970 4922
rect 2982 4870 3034 4922
rect 3046 4870 3098 4922
rect 3110 4870 3162 4922
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 6918 4870 6970 4922
rect 6982 4870 7034 4922
rect 7046 4870 7098 4922
rect 7110 4870 7162 4922
rect 7174 4870 7226 4922
rect 7238 4870 7290 4922
rect 10918 4870 10970 4922
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 11238 4870 11290 4922
rect 14918 4870 14970 4922
rect 14982 4870 15034 4922
rect 15046 4870 15098 4922
rect 15110 4870 15162 4922
rect 15174 4870 15226 4922
rect 15238 4870 15290 4922
rect 18918 4870 18970 4922
rect 18982 4870 19034 4922
rect 19046 4870 19098 4922
rect 19110 4870 19162 4922
rect 19174 4870 19226 4922
rect 19238 4870 19290 4922
rect 22918 4870 22970 4922
rect 22982 4870 23034 4922
rect 23046 4870 23098 4922
rect 23110 4870 23162 4922
rect 23174 4870 23226 4922
rect 23238 4870 23290 4922
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 6552 4768 6604 4820
rect 9220 4768 9272 4820
rect 5632 4700 5684 4752
rect 5264 4632 5316 4684
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 4436 4496 4488 4548
rect 5540 4564 5592 4616
rect 7564 4700 7616 4752
rect 5908 4564 5960 4616
rect 7932 4632 7984 4684
rect 11152 4700 11204 4752
rect 13820 4700 13872 4752
rect 14740 4811 14792 4820
rect 14740 4777 14749 4811
rect 14749 4777 14783 4811
rect 14783 4777 14792 4811
rect 14740 4768 14792 4777
rect 17224 4768 17276 4820
rect 19800 4768 19852 4820
rect 20352 4768 20404 4820
rect 20536 4768 20588 4820
rect 22100 4768 22152 4820
rect 18512 4743 18564 4752
rect 18512 4709 18521 4743
rect 18521 4709 18555 4743
rect 18555 4709 18564 4743
rect 18512 4700 18564 4709
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 10324 4632 10376 4684
rect 10692 4632 10744 4684
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 14924 4632 14976 4684
rect 6644 4539 6696 4548
rect 6644 4505 6653 4539
rect 6653 4505 6687 4539
rect 6687 4505 6696 4539
rect 6644 4496 6696 4505
rect 8300 4496 8352 4548
rect 9404 4496 9456 4548
rect 10784 4496 10836 4548
rect 2872 4428 2924 4480
rect 4528 4471 4580 4480
rect 4528 4437 4537 4471
rect 4537 4437 4571 4471
rect 4571 4437 4580 4471
rect 4528 4428 4580 4437
rect 7104 4428 7156 4480
rect 8392 4428 8444 4480
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 10232 4471 10284 4480
rect 10232 4437 10241 4471
rect 10241 4437 10275 4471
rect 10275 4437 10284 4471
rect 10232 4428 10284 4437
rect 10600 4428 10652 4480
rect 13636 4564 13688 4616
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 10968 4539 11020 4548
rect 10968 4505 10977 4539
rect 10977 4505 11011 4539
rect 11011 4505 11020 4539
rect 10968 4496 11020 4505
rect 11336 4428 11388 4480
rect 12992 4496 13044 4548
rect 13912 4496 13964 4548
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14648 4564 14700 4616
rect 16580 4564 16632 4616
rect 18328 4632 18380 4684
rect 16396 4496 16448 4548
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 19432 4564 19484 4616
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 17408 4496 17460 4548
rect 18788 4496 18840 4548
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 20812 4564 20864 4616
rect 20536 4496 20588 4548
rect 21916 4607 21968 4616
rect 21916 4573 21925 4607
rect 21925 4573 21959 4607
rect 21959 4573 21968 4607
rect 21916 4564 21968 4573
rect 22192 4607 22244 4616
rect 22192 4573 22201 4607
rect 22201 4573 22235 4607
rect 22235 4573 22244 4607
rect 22192 4564 22244 4573
rect 22652 4564 22704 4616
rect 24400 4564 24452 4616
rect 25228 4564 25280 4616
rect 24216 4496 24268 4548
rect 17868 4428 17920 4480
rect 20628 4428 20680 4480
rect 21088 4471 21140 4480
rect 21088 4437 21097 4471
rect 21097 4437 21131 4471
rect 21131 4437 21140 4471
rect 21088 4428 21140 4437
rect 22100 4428 22152 4480
rect 22560 4471 22612 4480
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 22560 4428 22612 4437
rect 23480 4428 23532 4480
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 3658 4326 3710 4378
rect 3722 4326 3774 4378
rect 3786 4326 3838 4378
rect 3850 4326 3902 4378
rect 3914 4326 3966 4378
rect 3978 4326 4030 4378
rect 7658 4326 7710 4378
rect 7722 4326 7774 4378
rect 7786 4326 7838 4378
rect 7850 4326 7902 4378
rect 7914 4326 7966 4378
rect 7978 4326 8030 4378
rect 11658 4326 11710 4378
rect 11722 4326 11774 4378
rect 11786 4326 11838 4378
rect 11850 4326 11902 4378
rect 11914 4326 11966 4378
rect 11978 4326 12030 4378
rect 15658 4326 15710 4378
rect 15722 4326 15774 4378
rect 15786 4326 15838 4378
rect 15850 4326 15902 4378
rect 15914 4326 15966 4378
rect 15978 4326 16030 4378
rect 19658 4326 19710 4378
rect 19722 4326 19774 4378
rect 19786 4326 19838 4378
rect 19850 4326 19902 4378
rect 19914 4326 19966 4378
rect 19978 4326 20030 4378
rect 23658 4326 23710 4378
rect 23722 4326 23774 4378
rect 23786 4326 23838 4378
rect 23850 4326 23902 4378
rect 23914 4326 23966 4378
rect 23978 4326 24030 4378
rect 5264 4224 5316 4276
rect 2872 4199 2924 4208
rect 2872 4165 2906 4199
rect 2906 4165 2924 4199
rect 2872 4156 2924 4165
rect 4528 4156 4580 4208
rect 1952 4088 2004 4140
rect 6368 4088 6420 4140
rect 8300 4267 8352 4276
rect 8300 4233 8309 4267
rect 8309 4233 8343 4267
rect 8343 4233 8352 4267
rect 8300 4224 8352 4233
rect 9128 4224 9180 4276
rect 10692 4224 10744 4276
rect 13176 4224 13228 4276
rect 13820 4224 13872 4276
rect 14096 4224 14148 4276
rect 16120 4267 16172 4276
rect 16120 4233 16129 4267
rect 16129 4233 16163 4267
rect 16163 4233 16172 4267
rect 16120 4224 16172 4233
rect 17316 4224 17368 4276
rect 17868 4224 17920 4276
rect 18144 4224 18196 4276
rect 20076 4267 20128 4276
rect 20076 4233 20085 4267
rect 20085 4233 20119 4267
rect 20119 4233 20128 4267
rect 20076 4224 20128 4233
rect 4436 3884 4488 3936
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 5632 3884 5684 3893
rect 8392 4088 8444 4140
rect 9496 4088 9548 4140
rect 10600 4131 10652 4140
rect 13268 4156 13320 4208
rect 16304 4156 16356 4208
rect 10600 4097 10618 4131
rect 10618 4097 10652 4131
rect 10600 4088 10652 4097
rect 11152 4131 11204 4140
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 13360 4088 13412 4140
rect 13728 4088 13780 4140
rect 6828 4020 6880 4072
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 11336 4020 11388 4072
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 16396 4088 16448 4140
rect 17408 4088 17460 4140
rect 17500 4088 17552 4140
rect 14924 4020 14976 4072
rect 16672 4020 16724 4072
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 18696 4156 18748 4208
rect 18604 4088 18656 4140
rect 19524 4131 19576 4140
rect 19524 4097 19533 4131
rect 19533 4097 19567 4131
rect 19567 4097 19576 4131
rect 19524 4088 19576 4097
rect 21088 4156 21140 4208
rect 22100 4199 22152 4208
rect 22100 4165 22109 4199
rect 22109 4165 22143 4199
rect 22143 4165 22152 4199
rect 22100 4156 22152 4165
rect 22560 4156 22612 4208
rect 19984 4088 20036 4140
rect 16212 3952 16264 4004
rect 18328 4020 18380 4072
rect 18512 3952 18564 4004
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 24216 4156 24268 4208
rect 24400 4156 24452 4208
rect 24952 4156 25004 4208
rect 25688 4088 25740 4140
rect 7104 3884 7156 3936
rect 10232 3884 10284 3936
rect 10600 3884 10652 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 15568 3884 15620 3936
rect 16120 3884 16172 3936
rect 17960 3884 18012 3936
rect 21456 3884 21508 3936
rect 22468 3884 22520 3936
rect 2918 3782 2970 3834
rect 2982 3782 3034 3834
rect 3046 3782 3098 3834
rect 3110 3782 3162 3834
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 6918 3782 6970 3834
rect 6982 3782 7034 3834
rect 7046 3782 7098 3834
rect 7110 3782 7162 3834
rect 7174 3782 7226 3834
rect 7238 3782 7290 3834
rect 10918 3782 10970 3834
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 11238 3782 11290 3834
rect 14918 3782 14970 3834
rect 14982 3782 15034 3834
rect 15046 3782 15098 3834
rect 15110 3782 15162 3834
rect 15174 3782 15226 3834
rect 15238 3782 15290 3834
rect 18918 3782 18970 3834
rect 18982 3782 19034 3834
rect 19046 3782 19098 3834
rect 19110 3782 19162 3834
rect 19174 3782 19226 3834
rect 19238 3782 19290 3834
rect 22918 3782 22970 3834
rect 22982 3782 23034 3834
rect 23046 3782 23098 3834
rect 23110 3782 23162 3834
rect 23174 3782 23226 3834
rect 23238 3782 23290 3834
rect 6644 3680 6696 3732
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 9496 3680 9548 3732
rect 10692 3612 10744 3664
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9220 3544 9272 3553
rect 12072 3544 12124 3596
rect 14188 3680 14240 3732
rect 13728 3544 13780 3596
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 16396 3723 16448 3732
rect 16396 3689 16405 3723
rect 16405 3689 16439 3723
rect 16439 3689 16448 3723
rect 16396 3680 16448 3689
rect 16764 3680 16816 3732
rect 17408 3680 17460 3732
rect 14740 3544 14792 3553
rect 18420 3544 18472 3596
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 6828 3519 6880 3528
rect 5172 3476 5224 3485
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9312 3476 9364 3528
rect 12440 3519 12492 3528
rect 12440 3485 12474 3519
rect 12474 3485 12492 3519
rect 5632 3408 5684 3460
rect 7196 3408 7248 3460
rect 8852 3408 8904 3460
rect 11336 3408 11388 3460
rect 12440 3476 12492 3485
rect 13268 3476 13320 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 14832 3476 14884 3528
rect 21916 3680 21968 3732
rect 24952 3723 25004 3732
rect 24952 3689 24961 3723
rect 24961 3689 24995 3723
rect 24995 3689 25004 3723
rect 24952 3680 25004 3689
rect 22744 3544 22796 3596
rect 4528 3383 4580 3392
rect 4528 3349 4537 3383
rect 4537 3349 4571 3383
rect 4571 3349 4580 3383
rect 4528 3340 4580 3349
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 12256 3340 12308 3392
rect 15384 3408 15436 3460
rect 16304 3408 16356 3460
rect 16212 3340 16264 3392
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 23020 3476 23072 3528
rect 22468 3408 22520 3460
rect 22744 3340 22796 3392
rect 24492 3383 24544 3392
rect 24492 3349 24501 3383
rect 24501 3349 24535 3383
rect 24535 3349 24544 3383
rect 24492 3340 24544 3349
rect 3658 3238 3710 3290
rect 3722 3238 3774 3290
rect 3786 3238 3838 3290
rect 3850 3238 3902 3290
rect 3914 3238 3966 3290
rect 3978 3238 4030 3290
rect 7658 3238 7710 3290
rect 7722 3238 7774 3290
rect 7786 3238 7838 3290
rect 7850 3238 7902 3290
rect 7914 3238 7966 3290
rect 7978 3238 8030 3290
rect 11658 3238 11710 3290
rect 11722 3238 11774 3290
rect 11786 3238 11838 3290
rect 11850 3238 11902 3290
rect 11914 3238 11966 3290
rect 11978 3238 12030 3290
rect 15658 3238 15710 3290
rect 15722 3238 15774 3290
rect 15786 3238 15838 3290
rect 15850 3238 15902 3290
rect 15914 3238 15966 3290
rect 15978 3238 16030 3290
rect 19658 3238 19710 3290
rect 19722 3238 19774 3290
rect 19786 3238 19838 3290
rect 19850 3238 19902 3290
rect 19914 3238 19966 3290
rect 19978 3238 20030 3290
rect 23658 3238 23710 3290
rect 23722 3238 23774 3290
rect 23786 3238 23838 3290
rect 23850 3238 23902 3290
rect 23914 3238 23966 3290
rect 23978 3238 24030 3290
rect 4712 3136 4764 3188
rect 5908 3136 5960 3188
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 6644 3136 6696 3188
rect 7196 3179 7248 3188
rect 7196 3145 7205 3179
rect 7205 3145 7239 3179
rect 7239 3145 7248 3179
rect 7196 3136 7248 3145
rect 5172 3068 5224 3120
rect 4528 3000 4580 3052
rect 6276 3000 6328 3052
rect 8208 3136 8260 3188
rect 9772 3136 9824 3188
rect 13268 3179 13320 3188
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 14188 3136 14240 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 16304 3179 16356 3188
rect 16304 3145 16313 3179
rect 16313 3145 16347 3179
rect 16347 3145 16356 3179
rect 16304 3136 16356 3145
rect 18328 3136 18380 3188
rect 22468 3136 22520 3188
rect 24308 3136 24360 3188
rect 9128 3068 9180 3120
rect 8392 3000 8444 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 12072 3068 12124 3120
rect 12256 3068 12308 3120
rect 13084 3068 13136 3120
rect 13728 3000 13780 3052
rect 7472 2932 7524 2984
rect 17960 3068 18012 3120
rect 18788 3068 18840 3120
rect 23480 3068 23532 3120
rect 15568 3043 15620 3052
rect 15568 3009 15577 3043
rect 15577 3009 15611 3043
rect 15611 3009 15620 3043
rect 15568 3000 15620 3009
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 22652 3000 22704 3052
rect 23020 3000 23072 3052
rect 24492 3000 24544 3052
rect 21456 2932 21508 2984
rect 4160 2796 4212 2848
rect 5908 2796 5960 2848
rect 14740 2796 14792 2848
rect 2918 2694 2970 2746
rect 2982 2694 3034 2746
rect 3046 2694 3098 2746
rect 3110 2694 3162 2746
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 6918 2694 6970 2746
rect 6982 2694 7034 2746
rect 7046 2694 7098 2746
rect 7110 2694 7162 2746
rect 7174 2694 7226 2746
rect 7238 2694 7290 2746
rect 10918 2694 10970 2746
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 11238 2694 11290 2746
rect 14918 2694 14970 2746
rect 14982 2694 15034 2746
rect 15046 2694 15098 2746
rect 15110 2694 15162 2746
rect 15174 2694 15226 2746
rect 15238 2694 15290 2746
rect 18918 2694 18970 2746
rect 18982 2694 19034 2746
rect 19046 2694 19098 2746
rect 19110 2694 19162 2746
rect 19174 2694 19226 2746
rect 19238 2694 19290 2746
rect 22918 2694 22970 2746
rect 22982 2694 23034 2746
rect 23046 2694 23098 2746
rect 23110 2694 23162 2746
rect 23174 2694 23226 2746
rect 23238 2694 23290 2746
rect 6276 2592 6328 2644
rect 8392 2524 8444 2576
rect 16212 2567 16264 2576
rect 16212 2533 16221 2567
rect 16221 2533 16255 2567
rect 16255 2533 16264 2567
rect 16212 2524 16264 2533
rect 13636 2456 13688 2508
rect 5816 2388 5868 2440
rect 8392 2388 8444 2440
rect 12808 2388 12860 2440
rect 16120 2388 16172 2440
rect 3658 2150 3710 2202
rect 3722 2150 3774 2202
rect 3786 2150 3838 2202
rect 3850 2150 3902 2202
rect 3914 2150 3966 2202
rect 3978 2150 4030 2202
rect 7658 2150 7710 2202
rect 7722 2150 7774 2202
rect 7786 2150 7838 2202
rect 7850 2150 7902 2202
rect 7914 2150 7966 2202
rect 7978 2150 8030 2202
rect 11658 2150 11710 2202
rect 11722 2150 11774 2202
rect 11786 2150 11838 2202
rect 11850 2150 11902 2202
rect 11914 2150 11966 2202
rect 11978 2150 12030 2202
rect 15658 2150 15710 2202
rect 15722 2150 15774 2202
rect 15786 2150 15838 2202
rect 15850 2150 15902 2202
rect 15914 2150 15966 2202
rect 15978 2150 16030 2202
rect 19658 2150 19710 2202
rect 19722 2150 19774 2202
rect 19786 2150 19838 2202
rect 19850 2150 19902 2202
rect 19914 2150 19966 2202
rect 19978 2150 20030 2202
rect 23658 2150 23710 2202
rect 23722 2150 23774 2202
rect 23786 2150 23838 2202
rect 23850 2150 23902 2202
rect 23914 2150 23966 2202
rect 23978 2150 24030 2202
<< metal2 >>
rect 9678 29458 9734 30115
rect 9678 29430 9812 29458
rect 9678 29315 9734 29430
rect 2916 27772 3292 27781
rect 2972 27770 2996 27772
rect 3052 27770 3076 27772
rect 3132 27770 3156 27772
rect 3212 27770 3236 27772
rect 2972 27718 2982 27770
rect 3226 27718 3236 27770
rect 2972 27716 2996 27718
rect 3052 27716 3076 27718
rect 3132 27716 3156 27718
rect 3212 27716 3236 27718
rect 2916 27707 3292 27716
rect 6916 27772 7292 27781
rect 6972 27770 6996 27772
rect 7052 27770 7076 27772
rect 7132 27770 7156 27772
rect 7212 27770 7236 27772
rect 6972 27718 6982 27770
rect 7226 27718 7236 27770
rect 6972 27716 6996 27718
rect 7052 27716 7076 27718
rect 7132 27716 7156 27718
rect 7212 27716 7236 27718
rect 6916 27707 7292 27716
rect 9784 27606 9812 29430
rect 10322 29315 10378 30115
rect 10966 29315 11022 30115
rect 11610 29458 11666 30115
rect 12254 29458 12310 30115
rect 14186 29458 14242 30115
rect 11610 29430 11744 29458
rect 11610 29315 11666 29430
rect 10336 27606 10364 29315
rect 10980 27962 11008 29315
rect 10796 27934 11008 27962
rect 10796 27606 10824 27934
rect 10916 27772 11292 27781
rect 10972 27770 10996 27772
rect 11052 27770 11076 27772
rect 11132 27770 11156 27772
rect 11212 27770 11236 27772
rect 10972 27718 10982 27770
rect 11226 27718 11236 27770
rect 10972 27716 10996 27718
rect 11052 27716 11076 27718
rect 11132 27716 11156 27718
rect 11212 27716 11236 27718
rect 10916 27707 11292 27716
rect 11716 27606 11744 29430
rect 12254 29430 12388 29458
rect 12254 29315 12310 29430
rect 12360 27606 12388 29430
rect 14186 29430 14320 29458
rect 14186 29315 14242 29430
rect 14292 27606 14320 29430
rect 17406 29315 17462 30115
rect 19982 29458 20038 30115
rect 19982 29430 20116 29458
rect 19982 29315 20038 29430
rect 14916 27772 15292 27781
rect 14972 27770 14996 27772
rect 15052 27770 15076 27772
rect 15132 27770 15156 27772
rect 15212 27770 15236 27772
rect 14972 27718 14982 27770
rect 15226 27718 15236 27770
rect 14972 27716 14996 27718
rect 15052 27716 15076 27718
rect 15132 27716 15156 27718
rect 15212 27716 15236 27718
rect 14916 27707 15292 27716
rect 17420 27606 17448 29315
rect 18916 27772 19292 27781
rect 18972 27770 18996 27772
rect 19052 27770 19076 27772
rect 19132 27770 19156 27772
rect 19212 27770 19236 27772
rect 18972 27718 18982 27770
rect 19226 27718 19236 27770
rect 18972 27716 18996 27718
rect 19052 27716 19076 27718
rect 19132 27716 19156 27718
rect 19212 27716 19236 27718
rect 18916 27707 19292 27716
rect 20088 27606 20116 29430
rect 20626 29315 20682 30115
rect 22558 29315 22614 30115
rect 24490 29315 24546 30115
rect 9772 27600 9824 27606
rect 9772 27542 9824 27548
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 10784 27600 10836 27606
rect 10784 27542 10836 27548
rect 11704 27600 11756 27606
rect 11704 27542 11756 27548
rect 12348 27600 12400 27606
rect 12348 27542 12400 27548
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 20640 27538 20668 29315
rect 20628 27532 20680 27538
rect 20628 27474 20680 27480
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 20536 27464 20588 27470
rect 20536 27406 20588 27412
rect 3656 27228 4032 27237
rect 3712 27226 3736 27228
rect 3792 27226 3816 27228
rect 3872 27226 3896 27228
rect 3952 27226 3976 27228
rect 3712 27174 3722 27226
rect 3966 27174 3976 27226
rect 3712 27172 3736 27174
rect 3792 27172 3816 27174
rect 3872 27172 3896 27174
rect 3952 27172 3976 27174
rect 3656 27163 4032 27172
rect 7656 27228 8032 27237
rect 7712 27226 7736 27228
rect 7792 27226 7816 27228
rect 7872 27226 7896 27228
rect 7952 27226 7976 27228
rect 7712 27174 7722 27226
rect 7966 27174 7976 27226
rect 7712 27172 7736 27174
rect 7792 27172 7816 27174
rect 7872 27172 7896 27174
rect 7952 27172 7976 27174
rect 7656 27163 8032 27172
rect 9784 27130 9812 27406
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 8760 26988 8812 26994
rect 8760 26930 8812 26936
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 2916 26684 3292 26693
rect 2972 26682 2996 26684
rect 3052 26682 3076 26684
rect 3132 26682 3156 26684
rect 3212 26682 3236 26684
rect 2972 26630 2982 26682
rect 3226 26630 3236 26682
rect 2972 26628 2996 26630
rect 3052 26628 3076 26630
rect 3132 26628 3156 26630
rect 3212 26628 3236 26630
rect 2916 26619 3292 26628
rect 3422 26480 3478 26489
rect 3422 26415 3478 26424
rect 2916 25596 3292 25605
rect 2972 25594 2996 25596
rect 3052 25594 3076 25596
rect 3132 25594 3156 25596
rect 3212 25594 3236 25596
rect 2972 25542 2982 25594
rect 3226 25542 3236 25594
rect 2972 25540 2996 25542
rect 3052 25540 3076 25542
rect 3132 25540 3156 25542
rect 3212 25540 3236 25542
rect 2916 25531 3292 25540
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 2148 24206 2176 24550
rect 2916 24508 3292 24517
rect 2972 24506 2996 24508
rect 3052 24506 3076 24508
rect 3132 24506 3156 24508
rect 3212 24506 3236 24508
rect 2972 24454 2982 24506
rect 3226 24454 3236 24506
rect 2972 24452 2996 24454
rect 3052 24452 3076 24454
rect 3132 24452 3156 24454
rect 3212 24452 3236 24454
rect 2916 24443 3292 24452
rect 1952 24200 2004 24206
rect 1952 24142 2004 24148
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 1964 23730 1992 24142
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1964 23186 1992 23666
rect 2916 23420 3292 23429
rect 2972 23418 2996 23420
rect 3052 23418 3076 23420
rect 3132 23418 3156 23420
rect 3212 23418 3236 23420
rect 2972 23366 2982 23418
rect 3226 23366 3236 23418
rect 2972 23364 2996 23366
rect 3052 23364 3076 23366
rect 3132 23364 3156 23366
rect 3212 23364 3236 23366
rect 2916 23355 3292 23364
rect 1952 23180 2004 23186
rect 1952 23122 2004 23128
rect 2320 23044 2372 23050
rect 2320 22986 2372 22992
rect 2332 22778 2360 22986
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3160 22778 3188 22918
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3344 22710 3372 24550
rect 3332 22704 3384 22710
rect 3332 22646 3384 22652
rect 2916 22332 3292 22341
rect 2972 22330 2996 22332
rect 3052 22330 3076 22332
rect 3132 22330 3156 22332
rect 3212 22330 3236 22332
rect 2972 22278 2982 22330
rect 3226 22278 3236 22330
rect 2972 22276 2996 22278
rect 3052 22276 3076 22278
rect 3132 22276 3156 22278
rect 3212 22276 3236 22278
rect 2916 22267 3292 22276
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2332 21554 2360 21830
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 1964 21010 1992 21490
rect 2700 21146 2728 21966
rect 2916 21244 3292 21253
rect 2972 21242 2996 21244
rect 3052 21242 3076 21244
rect 3132 21242 3156 21244
rect 3212 21242 3236 21244
rect 2972 21190 2982 21242
rect 3226 21190 3236 21242
rect 2972 21188 2996 21190
rect 3052 21188 3076 21190
rect 3132 21188 3156 21190
rect 3212 21188 3236 21190
rect 2916 21179 3292 21188
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 3344 20890 3372 22646
rect 2412 20868 2464 20874
rect 2412 20810 2464 20816
rect 3252 20862 3372 20890
rect 2424 20602 2452 20810
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 3252 20482 3280 20862
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3344 20602 3372 20742
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 3252 20454 3372 20482
rect 2916 20156 3292 20165
rect 2972 20154 2996 20156
rect 3052 20154 3076 20156
rect 3132 20154 3156 20156
rect 3212 20154 3236 20156
rect 2972 20102 2982 20154
rect 3226 20102 3236 20154
rect 2972 20100 2996 20102
rect 3052 20100 3076 20102
rect 3132 20100 3156 20102
rect 3212 20100 3236 20102
rect 2916 20091 3292 20100
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2424 19514 2452 19722
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1412 17785 1440 18158
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 2148 17678 2176 18566
rect 2516 18290 2544 19790
rect 3160 19514 3188 19790
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3344 19378 3372 20454
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 2916 19068 3292 19077
rect 2972 19066 2996 19068
rect 3052 19066 3076 19068
rect 3132 19066 3156 19068
rect 3212 19066 3236 19068
rect 2972 19014 2982 19066
rect 3226 19014 3236 19066
rect 2972 19012 2996 19014
rect 3052 19012 3076 19014
rect 3132 19012 3156 19014
rect 3212 19012 3236 19014
rect 2916 19003 3292 19012
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2792 18290 2820 18566
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 1504 17270 1532 17614
rect 2516 17270 2544 18226
rect 2916 17980 3292 17989
rect 2972 17978 2996 17980
rect 3052 17978 3076 17980
rect 3132 17978 3156 17980
rect 3212 17978 3236 17980
rect 2972 17926 2982 17978
rect 3226 17926 3236 17978
rect 2972 17924 2996 17926
rect 3052 17924 3076 17926
rect 3132 17924 3156 17926
rect 3212 17924 3236 17926
rect 2916 17915 3292 17924
rect 1492 17264 1544 17270
rect 1492 17206 1544 17212
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2240 16794 2268 17138
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2516 16574 2544 17206
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2792 16590 2820 17002
rect 2916 16892 3292 16901
rect 2972 16890 2996 16892
rect 3052 16890 3076 16892
rect 3132 16890 3156 16892
rect 3212 16890 3236 16892
rect 2972 16838 2982 16890
rect 3226 16838 3236 16890
rect 2972 16836 2996 16838
rect 3052 16836 3076 16838
rect 3132 16836 3156 16838
rect 3212 16836 3236 16838
rect 2916 16827 3292 16836
rect 2240 16546 2544 16574
rect 2780 16584 2832 16590
rect 2240 16182 2268 16546
rect 2780 16526 2832 16532
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2148 15162 2176 16050
rect 2240 15502 2268 16118
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2240 14958 2268 15438
rect 2792 15026 2820 15914
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 2916 15804 3292 15813
rect 2972 15802 2996 15804
rect 3052 15802 3076 15804
rect 3132 15802 3156 15804
rect 3212 15802 3236 15804
rect 2972 15750 2982 15802
rect 3226 15750 3236 15802
rect 2972 15748 2996 15750
rect 3052 15748 3076 15750
rect 3132 15748 3156 15750
rect 3212 15748 3236 15750
rect 2916 15739 3292 15748
rect 3344 15502 3372 15846
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3332 15088 3384 15094
rect 3436 15065 3464 26415
rect 4068 26376 4120 26382
rect 4068 26318 4120 26324
rect 4436 26376 4488 26382
rect 4436 26318 4488 26324
rect 3516 26240 3568 26246
rect 3516 26182 3568 26188
rect 3528 25838 3556 26182
rect 3656 26140 4032 26149
rect 3712 26138 3736 26140
rect 3792 26138 3816 26140
rect 3872 26138 3896 26140
rect 3952 26138 3976 26140
rect 3712 26086 3722 26138
rect 3966 26086 3976 26138
rect 3712 26084 3736 26086
rect 3792 26084 3816 26086
rect 3872 26084 3896 26086
rect 3952 26084 3976 26086
rect 3656 26075 4032 26084
rect 3516 25832 3568 25838
rect 3516 25774 3568 25780
rect 4080 25498 4108 26318
rect 4448 25974 4476 26318
rect 4816 26314 4844 26726
rect 4804 26308 4856 26314
rect 4804 26250 4856 26256
rect 5000 26042 5028 26930
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 6916 26684 7292 26693
rect 6972 26682 6996 26684
rect 7052 26682 7076 26684
rect 7132 26682 7156 26684
rect 7212 26682 7236 26684
rect 6972 26630 6982 26682
rect 7226 26630 7236 26682
rect 6972 26628 6996 26630
rect 7052 26628 7076 26630
rect 7132 26628 7156 26630
rect 7212 26628 7236 26630
rect 6916 26619 7292 26628
rect 5080 26580 5132 26586
rect 5080 26522 5132 26528
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 4436 25968 4488 25974
rect 4436 25910 4488 25916
rect 5092 25906 5120 26522
rect 5448 26444 5500 26450
rect 5448 26386 5500 26392
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 7196 26444 7248 26450
rect 7380 26444 7432 26450
rect 7248 26404 7380 26432
rect 7196 26386 7248 26392
rect 7380 26386 7432 26392
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 4988 25832 5040 25838
rect 4988 25774 5040 25780
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 5000 25362 5028 25774
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 3656 25052 4032 25061
rect 3712 25050 3736 25052
rect 3792 25050 3816 25052
rect 3872 25050 3896 25052
rect 3952 25050 3976 25052
rect 3712 24998 3722 25050
rect 3966 24998 3976 25050
rect 3712 24996 3736 24998
rect 3792 24996 3816 24998
rect 3872 24996 3896 24998
rect 3952 24996 3976 24998
rect 3656 24987 4032 24996
rect 3516 24812 3568 24818
rect 3516 24754 3568 24760
rect 3528 24070 3556 24754
rect 5000 24750 5028 25298
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3528 22642 3556 24006
rect 3656 23964 4032 23973
rect 3712 23962 3736 23964
rect 3792 23962 3816 23964
rect 3872 23962 3896 23964
rect 3952 23962 3976 23964
rect 3712 23910 3722 23962
rect 3966 23910 3976 23962
rect 3712 23908 3736 23910
rect 3792 23908 3816 23910
rect 3872 23908 3896 23910
rect 3952 23908 3976 23910
rect 3656 23899 4032 23908
rect 4080 23866 4108 24618
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4344 24132 4396 24138
rect 4344 24074 4396 24080
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4356 23730 4384 24074
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4632 23798 4660 24006
rect 4816 23866 4844 24142
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 5000 23798 5028 24686
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4988 23792 5040 23798
rect 4988 23734 5040 23740
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 3656 22876 4032 22885
rect 3712 22874 3736 22876
rect 3792 22874 3816 22876
rect 3872 22874 3896 22876
rect 3952 22874 3976 22876
rect 3712 22822 3722 22874
rect 3966 22822 3976 22874
rect 3712 22820 3736 22822
rect 3792 22820 3816 22822
rect 3872 22820 3896 22822
rect 3952 22820 3976 22822
rect 3656 22811 4032 22820
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 3988 22166 4016 22578
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3656 21788 4032 21797
rect 3712 21786 3736 21788
rect 3792 21786 3816 21788
rect 3872 21786 3896 21788
rect 3952 21786 3976 21788
rect 3712 21734 3722 21786
rect 3966 21734 3976 21786
rect 3712 21732 3736 21734
rect 3792 21732 3816 21734
rect 3872 21732 3896 21734
rect 3952 21732 3976 21734
rect 3656 21723 4032 21732
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3528 20534 3556 21286
rect 3988 20942 4016 21286
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3656 20700 4032 20709
rect 3712 20698 3736 20700
rect 3792 20698 3816 20700
rect 3872 20698 3896 20700
rect 3952 20698 3976 20700
rect 3712 20646 3722 20698
rect 3966 20646 3976 20698
rect 3712 20644 3736 20646
rect 3792 20644 3816 20646
rect 3872 20644 3896 20646
rect 3952 20644 3976 20646
rect 3656 20635 4032 20644
rect 3516 20528 3568 20534
rect 3516 20470 3568 20476
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3528 19310 3556 20334
rect 3988 20262 4016 20402
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3988 19854 4016 20198
rect 4080 19854 4108 23666
rect 4252 22160 4304 22166
rect 4252 22102 4304 22108
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4172 20330 4200 20742
rect 4264 20466 4292 22102
rect 4356 22098 4384 23666
rect 5092 23118 5120 25842
rect 5172 25696 5224 25702
rect 5172 25638 5224 25644
rect 5184 25226 5212 25638
rect 5460 25294 5488 26386
rect 6828 25968 6880 25974
rect 6828 25910 6880 25916
rect 6092 25900 6144 25906
rect 6092 25842 6144 25848
rect 5908 25696 5960 25702
rect 5908 25638 5960 25644
rect 5920 25294 5948 25638
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5172 25220 5224 25226
rect 5172 25162 5224 25168
rect 5080 23112 5132 23118
rect 5080 23054 5132 23060
rect 4620 22704 4672 22710
rect 4620 22646 4672 22652
rect 4436 22568 4488 22574
rect 4436 22510 4488 22516
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4356 21554 4384 22034
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4448 21146 4476 22510
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4160 20324 4212 20330
rect 4212 20284 4476 20312
rect 4160 20266 4212 20272
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3656 19612 4032 19621
rect 3712 19610 3736 19612
rect 3792 19610 3816 19612
rect 3872 19610 3896 19612
rect 3952 19610 3976 19612
rect 3712 19558 3722 19610
rect 3966 19558 3976 19610
rect 3712 19556 3736 19558
rect 3792 19556 3816 19558
rect 3872 19556 3896 19558
rect 3952 19556 3976 19558
rect 3656 19547 4032 19556
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3528 17882 3556 18702
rect 3656 18524 4032 18533
rect 3712 18522 3736 18524
rect 3792 18522 3816 18524
rect 3872 18522 3896 18524
rect 3952 18522 3976 18524
rect 3712 18470 3722 18522
rect 3966 18470 3976 18522
rect 3712 18468 3736 18470
rect 3792 18468 3816 18470
rect 3872 18468 3896 18470
rect 3952 18468 3976 18470
rect 3656 18459 4032 18468
rect 4080 18290 4108 19382
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4264 18630 4292 19314
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3656 17436 4032 17445
rect 3712 17434 3736 17436
rect 3792 17434 3816 17436
rect 3872 17434 3896 17436
rect 3952 17434 3976 17436
rect 3712 17382 3722 17434
rect 3966 17382 3976 17434
rect 3712 17380 3736 17382
rect 3792 17380 3816 17382
rect 3872 17380 3896 17382
rect 3952 17380 3976 17382
rect 3656 17371 4032 17380
rect 4172 17202 4200 18022
rect 4264 17610 4292 18566
rect 4356 18426 4384 18634
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4356 17134 4384 17682
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3332 15030 3384 15036
rect 3422 15056 3478 15065
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2916 14716 3292 14725
rect 2972 14714 2996 14716
rect 3052 14714 3076 14716
rect 3132 14714 3156 14716
rect 3212 14714 3236 14716
rect 2972 14662 2982 14714
rect 3226 14662 3236 14714
rect 2972 14660 2996 14662
rect 3052 14660 3076 14662
rect 3132 14660 3156 14662
rect 3212 14660 3236 14662
rect 2916 14651 3292 14660
rect 3344 14618 3372 15030
rect 3422 14991 3478 15000
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 2916 13628 3292 13637
rect 2972 13626 2996 13628
rect 3052 13626 3076 13628
rect 3132 13626 3156 13628
rect 3212 13626 3236 13628
rect 2972 13574 2982 13626
rect 3226 13574 3236 13626
rect 2972 13572 2996 13574
rect 3052 13572 3076 13574
rect 3132 13572 3156 13574
rect 3212 13572 3236 13574
rect 2916 13563 3292 13572
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2056 12986 2084 13262
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 846 12880 902 12889
rect 846 12815 848 12824
rect 900 12815 902 12824
rect 848 12786 900 12792
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11762 1624 12174
rect 2148 12170 2176 13126
rect 2792 12918 2820 13126
rect 2976 12986 3004 13262
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2332 12170 2360 12718
rect 2916 12540 3292 12549
rect 2972 12538 2996 12540
rect 3052 12538 3076 12540
rect 3132 12538 3156 12540
rect 3212 12538 3236 12540
rect 2972 12486 2982 12538
rect 3226 12486 3236 12538
rect 2972 12484 2996 12486
rect 3052 12484 3076 12486
rect 3132 12484 3156 12486
rect 3212 12484 3236 12486
rect 2916 12475 3292 12484
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2148 11354 2176 11698
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2608 11150 2636 11562
rect 2916 11452 3292 11461
rect 2972 11450 2996 11452
rect 3052 11450 3076 11452
rect 3132 11450 3156 11452
rect 3212 11450 3236 11452
rect 2972 11398 2982 11450
rect 3226 11398 3236 11450
rect 2972 11396 2996 11398
rect 3052 11396 3076 11398
rect 3132 11396 3156 11398
rect 3212 11396 3236 11398
rect 2916 11387 3292 11396
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 9625 1440 10542
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 10062 1532 10406
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 1492 10056 1544 10062
rect 2700 10033 2728 10066
rect 2792 10062 2820 10678
rect 2916 10364 3292 10373
rect 2972 10362 2996 10364
rect 3052 10362 3076 10364
rect 3132 10362 3156 10364
rect 3212 10362 3236 10364
rect 2972 10310 2982 10362
rect 3226 10310 3236 10362
rect 2972 10308 2996 10310
rect 3052 10308 3076 10310
rect 3132 10308 3156 10310
rect 3212 10308 3236 10310
rect 2916 10299 3292 10308
rect 3344 10266 3372 11630
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 2780 10056 2832 10062
rect 1492 9998 1544 10004
rect 2686 10024 2742 10033
rect 2780 9998 2832 10004
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 2686 9959 2742 9968
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 1398 9616 1454 9625
rect 1872 9586 1900 9862
rect 1398 9551 1454 9560
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1504 8974 1532 9454
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1688 8906 1716 9318
rect 2700 9178 2728 9522
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2792 8974 2820 9862
rect 3344 9722 3372 9998
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 2916 9276 3292 9285
rect 2972 9274 2996 9276
rect 3052 9274 3076 9276
rect 3132 9274 3156 9276
rect 3212 9274 3236 9276
rect 2972 9222 2982 9274
rect 3226 9222 3236 9274
rect 2972 9220 2996 9222
rect 3052 9220 3076 9222
rect 3132 9220 3156 9222
rect 3212 9220 3236 9222
rect 2916 9211 3292 9220
rect 3436 9110 3464 10678
rect 3528 10033 3556 17002
rect 4448 16998 4476 20284
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 3656 16348 4032 16357
rect 3712 16346 3736 16348
rect 3792 16346 3816 16348
rect 3872 16346 3896 16348
rect 3952 16346 3976 16348
rect 3712 16294 3722 16346
rect 3966 16294 3976 16346
rect 3712 16292 3736 16294
rect 3792 16292 3816 16294
rect 3872 16292 3896 16294
rect 3952 16292 3976 16294
rect 3656 16283 4032 16292
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3804 15706 3832 16050
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3656 15260 4032 15269
rect 3712 15258 3736 15260
rect 3792 15258 3816 15260
rect 3872 15258 3896 15260
rect 3952 15258 3976 15260
rect 3712 15206 3722 15258
rect 3966 15206 3976 15258
rect 3712 15204 3736 15206
rect 3792 15204 3816 15206
rect 3872 15204 3896 15206
rect 3952 15204 3976 15206
rect 3656 15195 4032 15204
rect 4172 15094 4200 15914
rect 4264 15706 4292 16526
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4356 15162 4384 16526
rect 4448 15366 4476 16934
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3656 14172 4032 14181
rect 3712 14170 3736 14172
rect 3792 14170 3816 14172
rect 3872 14170 3896 14172
rect 3952 14170 3976 14172
rect 3712 14118 3722 14170
rect 3966 14118 3976 14170
rect 3712 14116 3736 14118
rect 3792 14116 3816 14118
rect 3872 14116 3896 14118
rect 3952 14116 3976 14118
rect 3656 14107 4032 14116
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3656 13084 4032 13093
rect 3712 13082 3736 13084
rect 3792 13082 3816 13084
rect 3872 13082 3896 13084
rect 3952 13082 3976 13084
rect 3712 13030 3722 13082
rect 3966 13030 3976 13082
rect 3712 13028 3736 13030
rect 3792 13028 3816 13030
rect 3872 13028 3896 13030
rect 3952 13028 3976 13030
rect 3656 13019 4032 13028
rect 4080 12646 4108 13330
rect 4172 13274 4200 15030
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4356 14414 4384 14758
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4172 13246 4292 13274
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12238 4108 12582
rect 4172 12442 4200 13126
rect 4264 12764 4292 13246
rect 4344 12776 4396 12782
rect 4264 12736 4344 12764
rect 4344 12718 4396 12724
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3656 11996 4032 12005
rect 3712 11994 3736 11996
rect 3792 11994 3816 11996
rect 3872 11994 3896 11996
rect 3952 11994 3976 11996
rect 3712 11942 3722 11994
rect 3966 11942 3976 11994
rect 3712 11940 3736 11942
rect 3792 11940 3816 11942
rect 3872 11940 3896 11942
rect 3952 11940 3976 11942
rect 3656 11931 4032 11940
rect 3700 11688 3752 11694
rect 3698 11656 3700 11665
rect 3752 11656 3754 11665
rect 3698 11591 3754 11600
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 3656 10908 4032 10917
rect 3712 10906 3736 10908
rect 3792 10906 3816 10908
rect 3872 10906 3896 10908
rect 3952 10906 3976 10908
rect 3712 10854 3722 10906
rect 3966 10854 3976 10906
rect 3712 10852 3736 10854
rect 3792 10852 3816 10854
rect 3872 10852 3896 10854
rect 3952 10852 3976 10854
rect 3656 10843 4032 10852
rect 4172 10674 4200 10950
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3804 10062 3832 10610
rect 4448 10198 4476 13330
rect 4540 13326 4568 22374
rect 4632 21962 4660 22646
rect 5184 22030 5212 25162
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5276 24138 5304 24550
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 5368 23322 5396 24754
rect 5460 24206 5488 25230
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5724 23588 5776 23594
rect 5724 23530 5776 23536
rect 5356 23316 5408 23322
rect 5356 23258 5408 23264
rect 5540 23248 5592 23254
rect 5460 23196 5540 23202
rect 5460 23190 5592 23196
rect 5460 23174 5580 23190
rect 5736 23186 5764 23530
rect 5920 23186 5948 25094
rect 6104 24954 6132 25842
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 6472 24954 6500 25094
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 6564 24886 6592 25094
rect 6552 24880 6604 24886
rect 6552 24822 6604 24828
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 6012 23186 6040 23462
rect 5724 23180 5776 23186
rect 5460 23118 5488 23174
rect 5908 23180 5960 23186
rect 5724 23122 5776 23128
rect 5828 23140 5908 23168
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5264 23044 5316 23050
rect 5264 22986 5316 22992
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4632 19258 4660 21898
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 21622 4752 21830
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 4908 20602 4936 21966
rect 4896 20596 4948 20602
rect 5276 20584 5304 22986
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 5368 22137 5396 22918
rect 5354 22128 5410 22137
rect 5354 22063 5410 22072
rect 5460 21962 5488 23054
rect 5448 21956 5500 21962
rect 5448 21898 5500 21904
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 4896 20538 4948 20544
rect 5184 20556 5304 20584
rect 5184 20058 5212 20556
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4724 19446 4752 19790
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4632 19230 4752 19258
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4632 16590 4660 17206
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4724 16402 4752 19230
rect 4816 18766 4844 19654
rect 5276 19417 5304 20402
rect 5262 19408 5318 19417
rect 5262 19343 5318 19352
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4908 17678 4936 18702
rect 5000 18698 5028 18906
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4816 17202 4844 17478
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4632 16374 4752 16402
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4632 12434 4660 16374
rect 4816 16250 4844 17138
rect 5000 16658 5028 18634
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4724 15502 4752 16118
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4724 12889 4752 15438
rect 4816 14958 4844 16186
rect 5000 15502 5028 16458
rect 5092 15570 5120 18770
rect 5264 18760 5316 18766
rect 5184 18708 5264 18714
rect 5184 18702 5316 18708
rect 5184 18686 5304 18702
rect 5184 18086 5212 18686
rect 5368 18426 5396 21558
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5552 20618 5580 20810
rect 5460 20590 5580 20618
rect 5644 20602 5672 21286
rect 5736 20942 5764 21286
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5828 20806 5856 23140
rect 5908 23122 5960 23128
rect 6000 23180 6052 23186
rect 6000 23122 6052 23128
rect 6288 23118 6316 24006
rect 6564 23118 6592 24822
rect 6840 23866 6868 25910
rect 7024 25906 7052 26386
rect 7104 26240 7156 26246
rect 7104 26182 7156 26188
rect 7116 25974 7144 26182
rect 7104 25968 7156 25974
rect 7104 25910 7156 25916
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 6916 25596 7292 25605
rect 6972 25594 6996 25596
rect 7052 25594 7076 25596
rect 7132 25594 7156 25596
rect 7212 25594 7236 25596
rect 6972 25542 6982 25594
rect 7226 25542 7236 25594
rect 6972 25540 6996 25542
rect 7052 25540 7076 25542
rect 7132 25540 7156 25542
rect 7212 25540 7236 25542
rect 6916 25531 7292 25540
rect 7392 25362 7420 26386
rect 7668 26382 7696 26726
rect 7656 26376 7708 26382
rect 7656 26318 7708 26324
rect 7656 26140 8032 26149
rect 7712 26138 7736 26140
rect 7792 26138 7816 26140
rect 7872 26138 7896 26140
rect 7952 26138 7976 26140
rect 7712 26086 7722 26138
rect 7966 26086 7976 26138
rect 7712 26084 7736 26086
rect 7792 26084 7816 26086
rect 7872 26084 7896 26086
rect 7952 26084 7976 26086
rect 7656 26075 8032 26084
rect 7380 25356 7432 25362
rect 7380 25298 7432 25304
rect 7656 25052 8032 25061
rect 7712 25050 7736 25052
rect 7792 25050 7816 25052
rect 7872 25050 7896 25052
rect 7952 25050 7976 25052
rect 7712 24998 7722 25050
rect 7966 24998 7976 25050
rect 7712 24996 7736 24998
rect 7792 24996 7816 24998
rect 7872 24996 7896 24998
rect 7952 24996 7976 24998
rect 7656 24987 8032 24996
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 6916 24508 7292 24517
rect 6972 24506 6996 24508
rect 7052 24506 7076 24508
rect 7132 24506 7156 24508
rect 7212 24506 7236 24508
rect 6972 24454 6982 24506
rect 7226 24454 7236 24506
rect 6972 24452 6996 24454
rect 7052 24452 7076 24454
rect 7132 24452 7156 24454
rect 7212 24452 7236 24454
rect 6916 24443 7292 24452
rect 7576 24138 7604 24686
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6840 23594 6868 23802
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 6828 23588 6880 23594
rect 6828 23530 6880 23536
rect 6916 23420 7292 23429
rect 6972 23418 6996 23420
rect 7052 23418 7076 23420
rect 7132 23418 7156 23420
rect 7212 23418 7236 23420
rect 6972 23366 6982 23418
rect 7226 23366 7236 23418
rect 6972 23364 6996 23366
rect 7052 23364 7076 23366
rect 7132 23364 7156 23366
rect 7212 23364 7236 23366
rect 6916 23355 7292 23364
rect 7392 23322 7420 23666
rect 7576 23662 7604 24074
rect 7656 23964 8032 23973
rect 7712 23962 7736 23964
rect 7792 23962 7816 23964
rect 7872 23962 7896 23964
rect 7952 23962 7976 23964
rect 7712 23910 7722 23962
rect 7966 23910 7976 23962
rect 7712 23908 7736 23910
rect 7792 23908 7816 23910
rect 7872 23908 7896 23910
rect 7952 23908 7976 23910
rect 7656 23899 8032 23908
rect 8404 23662 8432 26862
rect 8588 26450 8616 26862
rect 8772 26586 8800 26930
rect 9312 26920 9364 26926
rect 9312 26862 9364 26868
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 9036 26580 9088 26586
rect 9036 26522 9088 26528
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8588 26234 8616 26386
rect 8588 26206 8708 26234
rect 8680 24750 8708 26206
rect 9048 25906 9076 26522
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9232 25702 9260 26726
rect 9324 26246 9352 26862
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9324 26042 9352 26182
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 8864 24954 8892 25298
rect 9232 25294 9260 25638
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9140 24954 9168 25230
rect 8852 24948 8904 24954
rect 8852 24890 8904 24896
rect 9128 24948 9180 24954
rect 9128 24890 9180 24896
rect 9232 24834 9260 25230
rect 9416 24886 9444 26182
rect 9692 25770 9720 26794
rect 9784 26042 9812 27066
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9680 25764 9732 25770
rect 9680 25706 9732 25712
rect 9956 25764 10008 25770
rect 9956 25706 10008 25712
rect 9968 25294 9996 25706
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9140 24806 9260 24834
rect 9404 24880 9456 24886
rect 9404 24822 9456 24828
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 8944 24744 8996 24750
rect 8944 24686 8996 24692
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 8116 23656 8168 23662
rect 8116 23598 8168 23604
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 7484 23474 7512 23598
rect 7484 23446 7604 23474
rect 7380 23316 7432 23322
rect 7432 23276 7512 23304
rect 7380 23258 7432 23264
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 7392 23050 7420 23122
rect 7380 23044 7432 23050
rect 7380 22986 7432 22992
rect 6184 22976 6236 22982
rect 6184 22918 6236 22924
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5920 21554 5948 21830
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5632 20596 5684 20602
rect 5460 19417 5488 20590
rect 5632 20538 5684 20544
rect 5828 20534 5856 20742
rect 5816 20528 5868 20534
rect 5816 20470 5868 20476
rect 5446 19408 5502 19417
rect 5446 19343 5448 19352
rect 5500 19343 5502 19352
rect 5448 19314 5500 19320
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 16182 5212 18022
rect 5368 17678 5396 18362
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5172 16176 5224 16182
rect 5172 16118 5224 16124
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13326 4844 13670
rect 4908 13462 4936 14894
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 5000 13394 5028 15438
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4804 13320 4856 13326
rect 4856 13268 4936 13274
rect 4804 13262 4936 13268
rect 4816 13246 4936 13262
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4816 12986 4844 13126
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4710 12880 4766 12889
rect 4710 12815 4766 12824
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4540 12406 4660 12434
rect 4540 11762 4568 12406
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4632 11898 4660 12106
rect 4724 12102 4752 12718
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4816 11762 4844 12582
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4908 11506 4936 13246
rect 4816 11478 4936 11506
rect 4816 10606 4844 11478
rect 5000 10810 5028 13330
rect 5092 10826 5120 15506
rect 5184 15502 5212 15982
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5276 13734 5304 16390
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5262 12880 5318 12889
rect 5262 12815 5318 12824
rect 5276 12782 5304 12815
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5368 12594 5396 16526
rect 5460 12850 5488 17546
rect 5552 16266 5580 18566
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 17882 5672 18226
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 6012 16794 6040 21422
rect 6196 21350 6224 22918
rect 7484 22642 7512 23276
rect 7576 23050 7604 23446
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 6460 22568 6512 22574
rect 6460 22510 6512 22516
rect 6472 22098 6500 22510
rect 6916 22332 7292 22341
rect 6972 22330 6996 22332
rect 7052 22330 7076 22332
rect 7132 22330 7156 22332
rect 7212 22330 7236 22332
rect 6972 22278 6982 22330
rect 7226 22278 7236 22330
rect 6972 22276 6996 22278
rect 7052 22276 7076 22278
rect 7132 22276 7156 22278
rect 7212 22276 7236 22278
rect 6916 22267 7292 22276
rect 7392 22234 7420 22578
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 6460 22092 6512 22098
rect 6460 22034 6512 22040
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6380 20330 6408 21490
rect 6472 21010 6500 22034
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6656 21350 6684 21490
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6656 19938 6684 21286
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 6748 20602 6776 20810
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6656 19910 6776 19938
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6092 19712 6144 19718
rect 6092 19654 6144 19660
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5552 16238 5672 16266
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5552 15570 5580 16118
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5644 13326 5672 16238
rect 5920 16114 5948 16390
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5908 15428 5960 15434
rect 5908 15370 5960 15376
rect 5920 15162 5948 15370
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5184 12566 5396 12594
rect 5184 11014 5212 12566
rect 5354 12472 5410 12481
rect 5354 12407 5410 12416
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4988 10804 5040 10810
rect 5092 10798 5212 10826
rect 4988 10746 5040 10752
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 3792 10056 3844 10062
rect 3514 10024 3570 10033
rect 3792 9998 3844 10004
rect 3514 9959 3570 9968
rect 3976 9920 4028 9926
rect 4028 9880 4108 9908
rect 3976 9862 4028 9868
rect 3656 9820 4032 9829
rect 3712 9818 3736 9820
rect 3792 9818 3816 9820
rect 3872 9818 3896 9820
rect 3952 9818 3976 9820
rect 3712 9766 3722 9818
rect 3966 9766 3976 9818
rect 3712 9764 3736 9766
rect 3792 9764 3816 9766
rect 3872 9764 3896 9766
rect 3952 9764 3976 9766
rect 3656 9755 4032 9764
rect 4080 9586 4108 9880
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3528 9042 3556 9522
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 1676 8900 1728 8906
rect 1676 8842 1728 8848
rect 3656 8732 4032 8741
rect 3712 8730 3736 8732
rect 3792 8730 3816 8732
rect 3872 8730 3896 8732
rect 3952 8730 3976 8732
rect 3712 8678 3722 8730
rect 3966 8678 3976 8730
rect 3712 8676 3736 8678
rect 3792 8676 3816 8678
rect 3872 8676 3896 8678
rect 3952 8676 3976 8678
rect 3656 8667 4032 8676
rect 2916 8188 3292 8197
rect 2972 8186 2996 8188
rect 3052 8186 3076 8188
rect 3132 8186 3156 8188
rect 3212 8186 3236 8188
rect 2972 8134 2982 8186
rect 3226 8134 3236 8186
rect 2972 8132 2996 8134
rect 3052 8132 3076 8134
rect 3132 8132 3156 8134
rect 3212 8132 3236 8134
rect 2916 8123 3292 8132
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3656 7644 4032 7653
rect 3712 7642 3736 7644
rect 3792 7642 3816 7644
rect 3872 7642 3896 7644
rect 3952 7642 3976 7644
rect 3712 7590 3722 7642
rect 3966 7590 3976 7642
rect 3712 7588 3736 7590
rect 3792 7588 3816 7590
rect 3872 7588 3896 7590
rect 3952 7588 3976 7590
rect 3656 7579 4032 7588
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6186 1440 6734
rect 1688 6322 1716 7142
rect 1872 6798 1900 7210
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6390 1900 6598
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 1964 6322 1992 6734
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1400 6180 1452 6186
rect 1400 6122 1452 6128
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5710 1808 6054
rect 1964 5914 1992 6258
rect 2792 5914 2820 7482
rect 4080 7478 4108 7754
rect 3516 7472 3568 7478
rect 4068 7472 4120 7478
rect 3516 7414 3568 7420
rect 3606 7440 3662 7449
rect 2916 7100 3292 7109
rect 2972 7098 2996 7100
rect 3052 7098 3076 7100
rect 3132 7098 3156 7100
rect 3212 7098 3236 7100
rect 2972 7046 2982 7098
rect 3226 7046 3236 7098
rect 2972 7044 2996 7046
rect 3052 7044 3076 7046
rect 3132 7044 3156 7046
rect 3212 7044 3236 7046
rect 2916 7035 3292 7044
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6390 3372 6598
rect 3436 6458 3464 6734
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3528 6118 3556 7414
rect 4068 7414 4120 7420
rect 3606 7375 3662 7384
rect 3620 7342 3648 7375
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3656 6556 4032 6565
rect 3712 6554 3736 6556
rect 3792 6554 3816 6556
rect 3872 6554 3896 6556
rect 3952 6554 3976 6556
rect 3712 6502 3722 6554
rect 3966 6502 3976 6554
rect 3712 6500 3736 6502
rect 3792 6500 3816 6502
rect 3872 6500 3896 6502
rect 3952 6500 3976 6502
rect 3656 6491 4032 6500
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 2916 6012 3292 6021
rect 2972 6010 2996 6012
rect 3052 6010 3076 6012
rect 3132 6010 3156 6012
rect 3212 6010 3236 6012
rect 2972 5958 2982 6010
rect 3226 5958 3236 6010
rect 2972 5956 2996 5958
rect 3052 5956 3076 5958
rect 3132 5956 3156 5958
rect 3212 5956 3236 5958
rect 2916 5947 3292 5956
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1964 4146 1992 5850
rect 4080 5846 4108 6190
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3656 5468 4032 5477
rect 3712 5466 3736 5468
rect 3792 5466 3816 5468
rect 3872 5466 3896 5468
rect 3952 5466 3976 5468
rect 3712 5414 3722 5466
rect 3966 5414 3976 5466
rect 3712 5412 3736 5414
rect 3792 5412 3816 5414
rect 3872 5412 3896 5414
rect 3952 5412 3976 5414
rect 3656 5403 4032 5412
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 2916 4924 3292 4933
rect 2972 4922 2996 4924
rect 3052 4922 3076 4924
rect 3132 4922 3156 4924
rect 3212 4922 3236 4924
rect 2972 4870 2982 4922
rect 3226 4870 3236 4922
rect 2972 4868 2996 4870
rect 3052 4868 3076 4870
rect 3132 4868 3156 4870
rect 3212 4868 3236 4870
rect 2916 4859 3292 4868
rect 3988 4622 4016 4966
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4214 2912 4422
rect 3656 4380 4032 4389
rect 3712 4378 3736 4380
rect 3792 4378 3816 4380
rect 3872 4378 3896 4380
rect 3952 4378 3976 4380
rect 3712 4326 3722 4378
rect 3966 4326 3976 4378
rect 3712 4324 3736 4326
rect 3792 4324 3816 4326
rect 3872 4324 3896 4326
rect 3952 4324 3976 4326
rect 3656 4315 4032 4324
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2916 3836 3292 3845
rect 2972 3834 2996 3836
rect 3052 3834 3076 3836
rect 3132 3834 3156 3836
rect 3212 3834 3236 3836
rect 2972 3782 2982 3834
rect 3226 3782 3236 3834
rect 2972 3780 2996 3782
rect 3052 3780 3076 3782
rect 3132 3780 3156 3782
rect 3212 3780 3236 3782
rect 2916 3771 3292 3780
rect 3656 3292 4032 3301
rect 3712 3290 3736 3292
rect 3792 3290 3816 3292
rect 3872 3290 3896 3292
rect 3952 3290 3976 3292
rect 3712 3238 3722 3290
rect 3966 3238 3976 3290
rect 3712 3236 3736 3238
rect 3792 3236 3816 3238
rect 3872 3236 3896 3238
rect 3952 3236 3976 3238
rect 3656 3227 4032 3236
rect 4172 2854 4200 10134
rect 4540 9926 4568 10202
rect 5092 10062 5120 10610
rect 5184 10130 5212 10798
rect 5368 10674 5396 12407
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4540 7546 4568 9862
rect 5000 8974 5028 9862
rect 5092 9178 5120 9998
rect 5276 9994 5304 10610
rect 5460 10282 5488 12650
rect 5552 12442 5580 12854
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5540 12436 5592 12442
rect 5644 12434 5672 12718
rect 5644 12406 5856 12434
rect 5540 12378 5592 12384
rect 5552 12322 5580 12378
rect 5552 12294 5672 12322
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5368 10266 5488 10282
rect 5356 10260 5488 10266
rect 5408 10254 5488 10260
rect 5356 10202 5408 10208
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5276 9722 5304 9930
rect 5460 9926 5488 10134
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5368 9722 5396 9862
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5184 8566 5212 9522
rect 5172 8560 5224 8566
rect 5170 8528 5172 8537
rect 5224 8528 5226 8537
rect 5170 8463 5226 8472
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4540 7449 4568 7482
rect 4526 7440 4582 7449
rect 5460 7410 5488 9862
rect 5552 9654 5580 12174
rect 5644 11762 5672 12294
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5736 11642 5764 11698
rect 5644 11614 5764 11642
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5552 8974 5580 9590
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 4526 7375 4582 7384
rect 5448 7404 5500 7410
rect 4540 6322 4568 7375
rect 5448 7346 5500 7352
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4448 4554 4476 5170
rect 4632 5166 4660 7278
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5170 7032 5226 7041
rect 5170 6967 5172 6976
rect 5224 6967 5226 6976
rect 5172 6938 5224 6944
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 6458 4752 6598
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 5184 5166 5212 6938
rect 5276 6798 5304 7142
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6390 5396 6734
rect 5460 6458 5488 7346
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4622 4752 4966
rect 5276 4690 5304 5170
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4448 3942 4476 4490
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4540 4214 4568 4422
rect 5276 4282 5304 4626
rect 5552 4622 5580 7754
rect 5644 4758 5672 11614
rect 5828 10554 5856 12406
rect 5920 11898 5948 13262
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6012 12306 6040 12718
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 6104 11762 6132 19654
rect 6564 19514 6592 19722
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6460 19440 6512 19446
rect 6460 19382 6512 19388
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6196 12986 6224 13262
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 5828 10526 6224 10554
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 5920 9994 5948 10406
rect 6104 10266 6132 10406
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5736 7449 5764 7482
rect 5722 7440 5778 7449
rect 5722 7375 5778 7384
rect 5828 6746 5856 9930
rect 6012 9586 6040 10134
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5920 8430 5948 8910
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6196 7342 6224 10526
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 5828 6718 5948 6746
rect 5920 6662 5948 6718
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6012 4826 6040 5170
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4540 3058 4568 3334
rect 4724 3194 4752 3470
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5184 3126 5212 3470
rect 5644 3466 5672 3878
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5920 3194 5948 4558
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 5920 2854 5948 3130
rect 6288 3058 6316 14554
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12918 6408 13126
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6380 11898 6408 12106
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 10062 6408 11494
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 8906 6408 9862
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6472 8514 6500 19382
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6564 17814 6592 18770
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6656 17746 6684 19790
rect 6748 19718 6776 19910
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6840 18272 6868 21490
rect 6916 21244 7292 21253
rect 6972 21242 6996 21244
rect 7052 21242 7076 21244
rect 7132 21242 7156 21244
rect 7212 21242 7236 21244
rect 6972 21190 6982 21242
rect 7226 21190 7236 21242
rect 6972 21188 6996 21190
rect 7052 21188 7076 21190
rect 7132 21188 7156 21190
rect 7212 21188 7236 21190
rect 6916 21179 7292 21188
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7392 20602 7420 20742
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 6916 20156 7292 20165
rect 6972 20154 6996 20156
rect 7052 20154 7076 20156
rect 7132 20154 7156 20156
rect 7212 20154 7236 20156
rect 6972 20102 6982 20154
rect 7226 20102 7236 20154
rect 6972 20100 6996 20102
rect 7052 20100 7076 20102
rect 7132 20100 7156 20102
rect 7212 20100 7236 20102
rect 6916 20091 7292 20100
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7024 19446 7052 19994
rect 7392 19938 7420 20538
rect 7116 19910 7420 19938
rect 7116 19446 7144 19910
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 7208 19378 7236 19654
rect 7380 19440 7432 19446
rect 7380 19382 7432 19388
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 7392 19242 7420 19382
rect 7576 19242 7604 22986
rect 7656 22876 8032 22885
rect 7712 22874 7736 22876
rect 7792 22874 7816 22876
rect 7872 22874 7896 22876
rect 7952 22874 7976 22876
rect 7712 22822 7722 22874
rect 7966 22822 7976 22874
rect 7712 22820 7736 22822
rect 7792 22820 7816 22822
rect 7872 22820 7896 22822
rect 7952 22820 7976 22822
rect 7656 22811 8032 22820
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8036 22030 8064 22374
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 8128 21894 8156 23598
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 8588 22710 8616 23190
rect 8772 23118 8800 23462
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8208 22092 8260 22098
rect 8312 22094 8340 22646
rect 8680 22098 8708 23054
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8772 22166 8800 22578
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8760 22160 8812 22166
rect 8760 22102 8812 22108
rect 8312 22066 8524 22094
rect 8208 22034 8260 22040
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 7656 21788 8032 21797
rect 7712 21786 7736 21788
rect 7792 21786 7816 21788
rect 7872 21786 7896 21788
rect 7952 21786 7976 21788
rect 7712 21734 7722 21786
rect 7966 21734 7976 21786
rect 7712 21732 7736 21734
rect 7792 21732 7816 21734
rect 7872 21732 7896 21734
rect 7952 21732 7976 21734
rect 7656 21723 8032 21732
rect 8128 20856 8156 21830
rect 8220 21622 8248 22034
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 8220 21146 8248 21558
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8128 20828 8432 20856
rect 7656 20700 8032 20709
rect 7712 20698 7736 20700
rect 7792 20698 7816 20700
rect 7872 20698 7896 20700
rect 7952 20698 7976 20700
rect 7712 20646 7722 20698
rect 7966 20646 7976 20698
rect 7712 20644 7736 20646
rect 7792 20644 7816 20646
rect 7872 20644 7896 20646
rect 7952 20644 7976 20646
rect 7656 20635 8032 20644
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7668 20058 7696 20538
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 7656 19612 8032 19621
rect 7712 19610 7736 19612
rect 7792 19610 7816 19612
rect 7872 19610 7896 19612
rect 7952 19610 7976 19612
rect 7712 19558 7722 19610
rect 7966 19558 7976 19610
rect 7712 19556 7736 19558
rect 7792 19556 7816 19558
rect 7872 19556 7896 19558
rect 7952 19556 7976 19558
rect 7656 19547 8032 19556
rect 8128 19514 8156 19654
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8220 19378 8248 20470
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 6916 19068 7292 19077
rect 6972 19066 6996 19068
rect 7052 19066 7076 19068
rect 7132 19066 7156 19068
rect 7212 19066 7236 19068
rect 6972 19014 6982 19066
rect 7226 19014 7236 19066
rect 6972 19012 6996 19014
rect 7052 19012 7076 19014
rect 7132 19012 7156 19014
rect 7212 19012 7236 19014
rect 6916 19003 7292 19012
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6748 18244 6868 18272
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6656 16250 6684 17682
rect 6748 17270 6776 18244
rect 6932 18170 6960 18566
rect 7024 18426 7052 18566
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6840 18142 6960 18170
rect 6840 17762 6868 18142
rect 7116 18086 7144 18226
rect 7208 18086 7236 18702
rect 7484 18426 7512 18702
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 6916 17980 7292 17989
rect 6972 17978 6996 17980
rect 7052 17978 7076 17980
rect 7132 17978 7156 17980
rect 7212 17978 7236 17980
rect 6972 17926 6982 17978
rect 7226 17926 7236 17978
rect 6972 17924 6996 17926
rect 7052 17924 7076 17926
rect 7132 17924 7156 17926
rect 7212 17924 7236 17926
rect 6916 17915 7292 17924
rect 6840 17734 6960 17762
rect 6932 17678 6960 17734
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6916 16892 7292 16901
rect 6972 16890 6996 16892
rect 7052 16890 7076 16892
rect 7132 16890 7156 16892
rect 7212 16890 7236 16892
rect 6972 16838 6982 16890
rect 7226 16838 7236 16890
rect 6972 16836 6996 16838
rect 7052 16836 7076 16838
rect 7132 16836 7156 16838
rect 7212 16836 7236 16838
rect 6916 16827 7292 16836
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6840 15042 6868 16594
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7116 16250 7144 16526
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7300 16182 7328 16458
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 6916 15804 7292 15813
rect 6972 15802 6996 15804
rect 7052 15802 7076 15804
rect 7132 15802 7156 15804
rect 7212 15802 7236 15804
rect 6972 15750 6982 15802
rect 7226 15750 7236 15802
rect 6972 15748 6996 15750
rect 7052 15748 7076 15750
rect 7132 15748 7156 15750
rect 7212 15748 7236 15750
rect 6916 15739 7292 15748
rect 7392 15706 7420 16458
rect 7576 16454 7604 18634
rect 7656 18524 8032 18533
rect 7712 18522 7736 18524
rect 7792 18522 7816 18524
rect 7872 18522 7896 18524
rect 7952 18522 7976 18524
rect 7712 18470 7722 18522
rect 7966 18470 7976 18522
rect 7712 18468 7736 18470
rect 7792 18468 7816 18470
rect 7872 18468 7896 18470
rect 7952 18468 7976 18470
rect 7656 18459 8032 18468
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8036 17882 8064 18226
rect 8128 18086 8156 19246
rect 8220 18850 8248 19314
rect 8220 18822 8340 18850
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 8220 18290 8248 18634
rect 8312 18630 8340 18822
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18426 8340 18566
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8312 18170 8340 18362
rect 8220 18142 8340 18170
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 7656 17436 8032 17445
rect 7712 17434 7736 17436
rect 7792 17434 7816 17436
rect 7872 17434 7896 17436
rect 7952 17434 7976 17436
rect 7712 17382 7722 17434
rect 7966 17382 7976 17434
rect 7712 17380 7736 17382
rect 7792 17380 7816 17382
rect 7872 17380 7896 17382
rect 7952 17380 7976 17382
rect 7656 17371 8032 17380
rect 8220 16726 8248 18142
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7656 16348 8032 16357
rect 7712 16346 7736 16348
rect 7792 16346 7816 16348
rect 7872 16346 7896 16348
rect 7952 16346 7976 16348
rect 7712 16294 7722 16346
rect 7966 16294 7976 16346
rect 7712 16292 7736 16294
rect 7792 16292 7816 16294
rect 7872 16292 7896 16294
rect 7952 16292 7976 16294
rect 7656 16283 8032 16292
rect 8220 16250 8248 16662
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 6932 15162 6960 15642
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6748 15014 6868 15042
rect 7024 15026 7052 15302
rect 7116 15162 7144 15370
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7012 15020 7064 15026
rect 6748 14550 6776 15014
rect 7012 14962 7064 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 6840 14618 6868 14894
rect 6916 14716 7292 14725
rect 6972 14714 6996 14716
rect 7052 14714 7076 14716
rect 7132 14714 7156 14716
rect 7212 14714 7236 14716
rect 6972 14662 6982 14714
rect 7226 14662 7236 14714
rect 6972 14660 6996 14662
rect 7052 14660 7076 14662
rect 7132 14660 7156 14662
rect 7212 14660 7236 14662
rect 6916 14651 7292 14660
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7484 14550 7512 14894
rect 7576 14890 7604 16050
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15502 8156 15846
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 7656 15260 8032 15269
rect 7712 15258 7736 15260
rect 7792 15258 7816 15260
rect 7872 15258 7896 15260
rect 7952 15258 7976 15260
rect 7712 15206 7722 15258
rect 7966 15206 7976 15258
rect 7712 15204 7736 15206
rect 7792 15204 7816 15206
rect 7872 15204 7896 15206
rect 7952 15204 7976 15206
rect 7656 15195 8032 15204
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7760 14929 7788 14962
rect 7746 14920 7802 14929
rect 7564 14884 7616 14890
rect 7746 14855 7802 14864
rect 7564 14826 7616 14832
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 11762 6592 13126
rect 6748 12918 6776 14486
rect 7656 14172 8032 14181
rect 7712 14170 7736 14172
rect 7792 14170 7816 14172
rect 7872 14170 7896 14172
rect 7952 14170 7976 14172
rect 7712 14118 7722 14170
rect 7966 14118 7976 14170
rect 7712 14116 7736 14118
rect 7792 14116 7816 14118
rect 7872 14116 7896 14118
rect 7952 14116 7976 14118
rect 7656 14107 8032 14116
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 6916 13628 7292 13637
rect 6972 13626 6996 13628
rect 7052 13626 7076 13628
rect 7132 13626 7156 13628
rect 7212 13626 7236 13628
rect 6972 13574 6982 13626
rect 7226 13574 7236 13626
rect 6972 13572 6996 13574
rect 7052 13572 7076 13574
rect 7132 13572 7156 13574
rect 7212 13572 7236 13574
rect 6916 13563 7292 13572
rect 7392 13462 7420 13942
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 7104 13388 7156 13394
rect 6840 13348 7104 13376
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6748 10198 6776 10610
rect 6840 10248 6868 13348
rect 7104 13330 7156 13336
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12918 6960 13126
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 6916 12540 7292 12549
rect 6972 12538 6996 12540
rect 7052 12538 7076 12540
rect 7132 12538 7156 12540
rect 7212 12538 7236 12540
rect 6972 12486 6982 12538
rect 7226 12486 7236 12538
rect 6972 12484 6996 12486
rect 7052 12484 7076 12486
rect 7132 12484 7156 12486
rect 7212 12484 7236 12486
rect 6916 12475 7292 12484
rect 7392 12442 7420 12854
rect 7576 12714 7604 13466
rect 7656 13084 8032 13093
rect 7712 13082 7736 13084
rect 7792 13082 7816 13084
rect 7872 13082 7896 13084
rect 7952 13082 7976 13084
rect 7712 13030 7722 13082
rect 7966 13030 7976 13082
rect 7712 13028 7736 13030
rect 7792 13028 7816 13030
rect 7872 13028 7896 13030
rect 7952 13028 7976 13030
rect 7656 13019 8032 13028
rect 8128 12866 8156 15302
rect 8312 15178 8340 16050
rect 8220 15162 8340 15178
rect 8208 15156 8340 15162
rect 8260 15150 8340 15156
rect 8208 15098 8260 15104
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8220 14618 8248 14962
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8036 12850 8156 12866
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 8024 12844 8156 12850
rect 8076 12838 8156 12844
rect 8024 12786 8076 12792
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7380 12436 7432 12442
rect 7668 12434 7696 12786
rect 8312 12782 8340 13398
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 7380 12378 7432 12384
rect 7576 12406 7696 12434
rect 6916 11452 7292 11461
rect 6972 11450 6996 11452
rect 7052 11450 7076 11452
rect 7132 11450 7156 11452
rect 7212 11450 7236 11452
rect 6972 11398 6982 11450
rect 7226 11398 7236 11450
rect 6972 11396 6996 11398
rect 7052 11396 7076 11398
rect 7132 11396 7156 11398
rect 7212 11396 7236 11398
rect 6916 11387 7292 11396
rect 7576 10810 7604 12406
rect 7656 11996 8032 12005
rect 7712 11994 7736 11996
rect 7792 11994 7816 11996
rect 7872 11994 7896 11996
rect 7952 11994 7976 11996
rect 7712 11942 7722 11994
rect 7966 11942 7976 11994
rect 7712 11940 7736 11942
rect 7792 11940 7816 11942
rect 7872 11940 7896 11942
rect 7952 11940 7976 11942
rect 7656 11931 8032 11940
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7656 10908 8032 10917
rect 7712 10906 7736 10908
rect 7792 10906 7816 10908
rect 7872 10906 7896 10908
rect 7952 10906 7976 10908
rect 7712 10854 7722 10906
rect 7966 10854 7976 10906
rect 7712 10852 7736 10854
rect 7792 10852 7816 10854
rect 7872 10852 7896 10854
rect 7952 10852 7976 10854
rect 7656 10843 8032 10852
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7208 10538 7236 10610
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 6916 10364 7292 10373
rect 6972 10362 6996 10364
rect 7052 10362 7076 10364
rect 7132 10362 7156 10364
rect 7212 10362 7236 10364
rect 6972 10310 6982 10362
rect 7226 10310 7236 10362
rect 6972 10308 6996 10310
rect 7052 10308 7076 10310
rect 7132 10308 7156 10310
rect 7212 10308 7236 10310
rect 6916 10299 7292 10308
rect 6840 10220 7236 10248
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 7102 10160 7158 10169
rect 7208 10130 7236 10220
rect 7102 10095 7104 10104
rect 7156 10095 7158 10104
rect 7196 10124 7248 10130
rect 7104 10066 7156 10072
rect 7196 10066 7248 10072
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 7208 9674 7236 10066
rect 7392 9994 7420 10678
rect 8128 10674 8156 10950
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8114 10568 8170 10577
rect 7472 10532 7524 10538
rect 8114 10503 8170 10512
rect 7472 10474 7524 10480
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 6840 9160 6868 9658
rect 7208 9646 7328 9674
rect 7300 9466 7328 9646
rect 7392 9586 7420 9930
rect 7484 9654 7512 10474
rect 7562 10296 7618 10305
rect 7562 10231 7564 10240
rect 7616 10231 7618 10240
rect 7564 10202 7616 10208
rect 8128 10146 8156 10503
rect 8220 10266 8248 11086
rect 8312 10577 8340 12718
rect 8298 10568 8354 10577
rect 8298 10503 8354 10512
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8128 10118 8248 10146
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9722 7604 9998
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 7656 9820 8032 9829
rect 7712 9818 7736 9820
rect 7792 9818 7816 9820
rect 7872 9818 7896 9820
rect 7952 9818 7976 9820
rect 7712 9766 7722 9818
rect 7966 9766 7976 9818
rect 7712 9764 7736 9766
rect 7792 9764 7816 9766
rect 7872 9764 7896 9766
rect 7952 9764 7976 9766
rect 7656 9755 8032 9764
rect 8128 9722 8156 9862
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7300 9438 7420 9466
rect 6916 9276 7292 9285
rect 6972 9274 6996 9276
rect 7052 9274 7076 9276
rect 7132 9274 7156 9276
rect 7212 9274 7236 9276
rect 6972 9222 6982 9274
rect 7226 9222 7236 9274
rect 6972 9220 6996 9222
rect 7052 9220 7076 9222
rect 7132 9220 7156 9222
rect 7212 9220 7236 9222
rect 6916 9211 7292 9220
rect 6840 9132 6960 9160
rect 6472 8486 6592 8514
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6472 7886 6500 8366
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6472 6798 6500 7822
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6380 5574 6408 6734
rect 6472 6390 6500 6734
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6564 4826 6592 8486
rect 6932 8378 6960 9132
rect 7392 8650 7420 9438
rect 7484 9178 7512 9590
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7656 8732 8032 8741
rect 7712 8730 7736 8732
rect 7792 8730 7816 8732
rect 7872 8730 7896 8732
rect 7952 8730 7976 8732
rect 7712 8678 7722 8730
rect 7966 8678 7976 8730
rect 7712 8676 7736 8678
rect 7792 8676 7816 8678
rect 7872 8676 7896 8678
rect 7952 8676 7976 8678
rect 7656 8667 8032 8676
rect 7392 8622 7604 8650
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 6840 8350 6960 8378
rect 6840 7970 6868 8350
rect 6916 8188 7292 8197
rect 6972 8186 6996 8188
rect 7052 8186 7076 8188
rect 7132 8186 7156 8188
rect 7212 8186 7236 8188
rect 6972 8134 6982 8186
rect 7226 8134 7236 8186
rect 6972 8132 6996 8134
rect 7052 8132 7076 8134
rect 7132 8132 7156 8134
rect 7212 8132 7236 8134
rect 6916 8123 7292 8132
rect 6840 7942 6960 7970
rect 6932 7426 6960 7942
rect 7392 7546 7420 8434
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 7886 7512 8230
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7380 7540 7432 7546
rect 7576 7528 7604 8622
rect 8220 7818 8248 10118
rect 8312 10062 8340 10406
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8404 9926 8432 20828
rect 8496 18766 8524 22066
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8588 21690 8616 21966
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8588 19854 8616 20198
rect 8680 19922 8708 22034
rect 8772 20806 8800 22102
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8772 19446 8800 20742
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8772 18834 8800 19110
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8588 17882 8616 18158
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8496 15026 8524 15438
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8484 14884 8536 14890
rect 8772 14872 8800 14962
rect 8536 14844 8800 14872
rect 8484 14826 8536 14832
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8496 12306 8524 12718
rect 8588 12442 8616 12786
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8772 12238 8800 13126
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8496 10033 8524 10066
rect 8576 10056 8628 10062
rect 8482 10024 8538 10033
rect 8576 9998 8628 10004
rect 8482 9959 8538 9968
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7656 7644 8032 7653
rect 7712 7642 7736 7644
rect 7792 7642 7816 7644
rect 7872 7642 7896 7644
rect 7952 7642 7976 7644
rect 7712 7590 7722 7642
rect 7966 7590 7976 7642
rect 7712 7588 7736 7590
rect 7792 7588 7816 7590
rect 7872 7588 7896 7590
rect 7952 7588 7976 7590
rect 7656 7579 8032 7588
rect 8128 7546 8156 7686
rect 7380 7482 7432 7488
rect 7484 7500 7604 7528
rect 8116 7540 8168 7546
rect 6932 7398 7420 7426
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6748 6798 6776 7142
rect 6840 7002 6868 7278
rect 6916 7100 7292 7109
rect 6972 7098 6996 7100
rect 7052 7098 7076 7100
rect 7132 7098 7156 7100
rect 7212 7098 7236 7100
rect 6972 7046 6982 7098
rect 7226 7046 7236 7098
rect 6972 7044 6996 7046
rect 7052 7044 7076 7046
rect 7132 7044 7156 7046
rect 7212 7044 7236 7046
rect 6916 7035 7292 7044
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 5914 6684 6258
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6380 3194 6408 4082
rect 6656 3738 6684 4490
rect 6840 4078 6868 6326
rect 7392 6254 7420 7398
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 6916 6012 7292 6021
rect 6972 6010 6996 6012
rect 7052 6010 7076 6012
rect 7132 6010 7156 6012
rect 7212 6010 7236 6012
rect 6972 5958 6982 6010
rect 7226 5958 7236 6010
rect 6972 5956 6996 5958
rect 7052 5956 7076 5958
rect 7132 5956 7156 5958
rect 7212 5956 7236 5958
rect 6916 5947 7292 5956
rect 7484 5030 7512 7500
rect 8116 7482 8168 7488
rect 8312 7449 8340 9522
rect 7746 7440 7802 7449
rect 7564 7404 7616 7410
rect 8298 7440 8354 7449
rect 7746 7375 7802 7384
rect 8208 7404 8260 7410
rect 7564 7346 7616 7352
rect 7576 7002 7604 7346
rect 7760 7342 7788 7375
rect 8588 7410 8616 9998
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8298 7375 8354 7384
rect 8392 7404 8444 7410
rect 8208 7346 8260 7352
rect 8392 7346 8444 7352
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8036 7002 8064 7278
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 8220 6934 8248 7346
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 6934 8340 7210
rect 8404 6934 8432 7346
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8220 6798 8248 6870
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 7656 6556 8032 6565
rect 7712 6554 7736 6556
rect 7792 6554 7816 6556
rect 7872 6554 7896 6556
rect 7952 6554 7976 6556
rect 7712 6502 7722 6554
rect 7966 6502 7976 6554
rect 7712 6500 7736 6502
rect 7792 6500 7816 6502
rect 7872 6500 7896 6502
rect 7952 6500 7976 6502
rect 7656 6491 8032 6500
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7576 5642 7604 6054
rect 7852 5710 7880 6054
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 6916 4924 7292 4933
rect 6972 4922 6996 4924
rect 7052 4922 7076 4924
rect 7132 4922 7156 4924
rect 7212 4922 7236 4924
rect 6972 4870 6982 4922
rect 7226 4870 7236 4922
rect 6972 4868 6996 4870
rect 7052 4868 7076 4870
rect 7132 4868 7156 4870
rect 7212 4868 7236 4870
rect 6916 4859 7292 4868
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6656 3194 6684 3674
rect 6840 3534 6868 4014
rect 7116 3942 7144 4422
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6916 3836 7292 3845
rect 6972 3834 6996 3836
rect 7052 3834 7076 3836
rect 7132 3834 7156 3836
rect 7212 3834 7236 3836
rect 6972 3782 6982 3834
rect 7226 3782 7236 3834
rect 6972 3780 6996 3782
rect 7052 3780 7076 3782
rect 7132 3780 7156 3782
rect 7212 3780 7236 3782
rect 6916 3771 7292 3780
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7208 3194 7236 3402
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 2916 2748 3292 2757
rect 2972 2746 2996 2748
rect 3052 2746 3076 2748
rect 3132 2746 3156 2748
rect 3212 2746 3236 2748
rect 2972 2694 2982 2746
rect 3226 2694 3236 2746
rect 2972 2692 2996 2694
rect 3052 2692 3076 2694
rect 3132 2692 3156 2694
rect 3212 2692 3236 2694
rect 2916 2683 3292 2692
rect 6288 2650 6316 2994
rect 7484 2990 7512 4966
rect 7576 4758 7604 5578
rect 8128 5574 8156 6598
rect 8496 6458 8524 7346
rect 8680 6798 8708 9862
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8498 8800 8774
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8680 6390 8708 6734
rect 8772 6390 8800 7142
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8680 5914 8708 6326
rect 8864 6118 8892 22374
rect 8956 21554 8984 24686
rect 9140 22438 9168 24806
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9508 22778 9536 23054
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9692 22658 9720 23122
rect 9600 22642 9720 22658
rect 9588 22636 9720 22642
rect 9640 22630 9720 22636
rect 9588 22578 9640 22584
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 22234 9168 22374
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 9508 21894 9536 22510
rect 9968 22438 9996 25230
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9508 21690 9536 21830
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9140 18970 9168 19110
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9324 18766 9352 19110
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8956 17066 8984 17546
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 8956 15094 8984 16118
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9048 15434 9076 15846
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 9140 15201 9168 18634
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9211 18352 9263 18358
rect 9324 18340 9352 18566
rect 9263 18312 9352 18340
rect 9211 18294 9263 18300
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9126 15192 9182 15201
rect 9126 15127 9182 15136
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8956 13462 8984 15030
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9048 14929 9076 14962
rect 9034 14920 9090 14929
rect 9034 14855 9090 14864
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 9232 12918 9260 17818
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9416 12434 9444 21422
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9508 17882 9536 18702
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9508 13462 9536 17002
rect 9600 15706 9628 20878
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9692 18873 9720 19178
rect 9678 18864 9734 18873
rect 9678 18799 9734 18808
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 18358 9720 18702
rect 9784 18426 9812 20878
rect 10060 20398 10088 21558
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9968 18970 9996 19314
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9692 17202 9720 18294
rect 9784 17678 9812 18362
rect 9876 18170 9904 18906
rect 9876 18142 9996 18170
rect 9968 18086 9996 18142
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 16794 9720 17138
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9692 16658 9720 16730
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9692 15502 9720 16594
rect 9784 16046 9812 17478
rect 10060 16182 10088 17682
rect 10048 16176 10100 16182
rect 9968 16124 10048 16130
rect 9968 16118 10100 16124
rect 9968 16102 10088 16118
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9784 14822 9812 15982
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9876 15162 9904 15370
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9600 13394 9628 14418
rect 9784 14346 9812 14758
rect 9876 14414 9904 15098
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9232 12406 9444 12434
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8956 10742 8984 12242
rect 9126 11792 9182 11801
rect 9126 11727 9182 11736
rect 9140 11150 9168 11727
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8956 10130 8984 10678
rect 9034 10160 9090 10169
rect 8944 10124 8996 10130
rect 9034 10095 9090 10104
rect 8944 10066 8996 10072
rect 8956 9586 8984 10066
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 8498 8984 9522
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 7954 8984 8434
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 9048 7834 9076 10095
rect 9232 9518 9260 12406
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9416 11898 9444 12106
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11150 9444 11630
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9324 10470 9352 11086
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10674 9628 10950
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9042 9260 9454
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 8956 7806 9076 7834
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8956 5930 8984 7806
rect 9140 7546 9168 7822
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9416 6458 9444 10610
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9508 10305 9536 10474
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9494 10296 9550 10305
rect 9494 10231 9550 10240
rect 9600 10033 9628 10406
rect 9586 10024 9642 10033
rect 9586 9959 9642 9968
rect 9692 9110 9720 11834
rect 9784 10656 9812 13806
rect 9968 13394 9996 16102
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9876 12646 9904 13194
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9968 12434 9996 12786
rect 9876 12406 9996 12434
rect 9876 11898 9904 12406
rect 10060 12374 10088 15982
rect 10048 12368 10100 12374
rect 9968 12316 10048 12322
rect 9968 12310 10100 12316
rect 9968 12294 10088 12310
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9864 10668 9916 10674
rect 9784 10628 9864 10656
rect 9864 10610 9916 10616
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9508 6322 9536 8910
rect 9692 6662 9720 9046
rect 9968 7206 9996 12294
rect 10046 10840 10102 10849
rect 10152 10810 10180 22918
rect 10244 21146 10272 26930
rect 10612 26926 10640 27406
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10784 27056 10836 27062
rect 11072 27010 11100 27066
rect 10784 26998 10836 27004
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10428 26042 10456 26386
rect 10520 26314 10548 26726
rect 10508 26308 10560 26314
rect 10508 26250 10560 26256
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10428 25226 10456 25978
rect 10704 25702 10732 26930
rect 10796 26858 10824 26998
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10980 26982 11100 27010
rect 10888 26897 10916 26930
rect 10874 26888 10930 26897
rect 10784 26852 10836 26858
rect 10874 26823 10930 26832
rect 10784 26794 10836 26800
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10508 25220 10560 25226
rect 10508 25162 10560 25168
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 24818 10364 25094
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10336 23118 10364 24618
rect 10428 23186 10456 25162
rect 10520 24954 10548 25162
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10796 24834 10824 26794
rect 10980 26790 11008 26982
rect 10968 26784 11020 26790
rect 10968 26726 11020 26732
rect 11336 26784 11388 26790
rect 11336 26726 11388 26732
rect 10916 26684 11292 26693
rect 10972 26682 10996 26684
rect 11052 26682 11076 26684
rect 11132 26682 11156 26684
rect 11212 26682 11236 26684
rect 10972 26630 10982 26682
rect 11226 26630 11236 26682
rect 10972 26628 10996 26630
rect 11052 26628 11076 26630
rect 11132 26628 11156 26630
rect 11212 26628 11236 26630
rect 10916 26619 11292 26628
rect 11348 26234 11376 26726
rect 11164 26206 11376 26234
rect 11164 25974 11192 26206
rect 11152 25968 11204 25974
rect 11152 25910 11204 25916
rect 10916 25596 11292 25605
rect 10972 25594 10996 25596
rect 11052 25594 11076 25596
rect 11132 25594 11156 25596
rect 11212 25594 11236 25596
rect 10972 25542 10982 25594
rect 11226 25542 11236 25594
rect 10972 25540 10996 25542
rect 11052 25540 11076 25542
rect 11132 25540 11156 25542
rect 11212 25540 11236 25542
rect 10916 25531 11292 25540
rect 10704 24818 10824 24834
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10692 24812 10824 24818
rect 10744 24806 10824 24812
rect 10692 24754 10744 24760
rect 10416 23180 10468 23186
rect 10416 23122 10468 23128
rect 10324 23112 10376 23118
rect 10376 23060 10456 23066
rect 10324 23054 10456 23060
rect 10336 23038 10456 23054
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10336 22574 10364 22918
rect 10428 22574 10456 23038
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10336 19718 10364 20402
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10336 19514 10364 19654
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10414 19408 10470 19417
rect 10414 19343 10416 19352
rect 10468 19343 10470 19352
rect 10416 19314 10468 19320
rect 10232 19304 10284 19310
rect 10230 19272 10232 19281
rect 10284 19272 10286 19281
rect 10230 19207 10286 19216
rect 10322 18864 10378 18873
rect 10322 18799 10378 18808
rect 10336 17882 10364 18799
rect 10428 18290 10456 19314
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10428 18193 10456 18226
rect 10414 18184 10470 18193
rect 10414 18119 10470 18128
rect 10520 17898 10548 24754
rect 10704 24682 10732 24754
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10916 24508 11292 24517
rect 10972 24506 10996 24508
rect 11052 24506 11076 24508
rect 11132 24506 11156 24508
rect 11212 24506 11236 24508
rect 10972 24454 10982 24506
rect 11226 24454 11236 24506
rect 10972 24452 10996 24454
rect 11052 24452 11076 24454
rect 11132 24452 11156 24454
rect 11212 24452 11236 24454
rect 10916 24443 11292 24452
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 10916 23420 11292 23429
rect 10972 23418 10996 23420
rect 11052 23418 11076 23420
rect 11132 23418 11156 23420
rect 11212 23418 11236 23420
rect 10972 23366 10982 23418
rect 11226 23366 11236 23418
rect 10972 23364 10996 23366
rect 11052 23364 11076 23366
rect 11132 23364 11156 23366
rect 11212 23364 11236 23366
rect 10916 23355 11292 23364
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10888 23089 10916 23258
rect 10874 23080 10930 23089
rect 10692 23044 10744 23050
rect 10874 23015 10930 23024
rect 10692 22986 10744 22992
rect 10704 22778 10732 22986
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 11348 22710 11376 23462
rect 11440 22982 11468 27338
rect 11532 25158 11560 27406
rect 11656 27228 12032 27237
rect 11712 27226 11736 27228
rect 11792 27226 11816 27228
rect 11872 27226 11896 27228
rect 11952 27226 11976 27228
rect 11712 27174 11722 27226
rect 11966 27174 11976 27226
rect 11712 27172 11736 27174
rect 11792 27172 11816 27174
rect 11872 27172 11896 27174
rect 11952 27172 11976 27174
rect 11656 27163 12032 27172
rect 11888 26920 11940 26926
rect 11888 26862 11940 26868
rect 11900 26586 11928 26862
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11656 26140 12032 26149
rect 11712 26138 11736 26140
rect 11792 26138 11816 26140
rect 11872 26138 11896 26140
rect 11952 26138 11976 26140
rect 11712 26086 11722 26138
rect 11966 26086 11976 26138
rect 11712 26084 11736 26086
rect 11792 26084 11816 26086
rect 11872 26084 11896 26086
rect 11952 26084 11976 26086
rect 11656 26075 12032 26084
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11532 24750 11560 25094
rect 11656 25052 12032 25061
rect 11712 25050 11736 25052
rect 11792 25050 11816 25052
rect 11872 25050 11896 25052
rect 11952 25050 11976 25052
rect 11712 24998 11722 25050
rect 11966 24998 11976 25050
rect 11712 24996 11736 24998
rect 11792 24996 11816 24998
rect 11872 24996 11896 24998
rect 11952 24996 11976 24998
rect 11656 24987 12032 24996
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11656 23964 12032 23973
rect 11712 23962 11736 23964
rect 11792 23962 11816 23964
rect 11872 23962 11896 23964
rect 11952 23962 11976 23964
rect 11712 23910 11722 23962
rect 11966 23910 11976 23962
rect 11712 23908 11736 23910
rect 11792 23908 11816 23910
rect 11872 23908 11896 23910
rect 11952 23908 11976 23910
rect 11656 23899 12032 23908
rect 12176 23322 12204 27406
rect 12532 27056 12584 27062
rect 12532 26998 12584 27004
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12268 25906 12296 26318
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 12268 25294 12296 25842
rect 12348 25356 12400 25362
rect 12348 25298 12400 25304
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12268 23730 12296 25230
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12268 23322 12296 23666
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11440 22574 11468 22918
rect 11656 22876 12032 22885
rect 11712 22874 11736 22876
rect 11792 22874 11816 22876
rect 11872 22874 11896 22876
rect 11952 22874 11976 22876
rect 11712 22822 11722 22874
rect 11966 22822 11976 22874
rect 11712 22820 11736 22822
rect 11792 22820 11816 22822
rect 11872 22820 11896 22822
rect 11952 22820 11976 22822
rect 11656 22811 12032 22820
rect 12176 22778 12204 23258
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12268 22710 12296 23122
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 10916 22332 11292 22341
rect 10972 22330 10996 22332
rect 11052 22330 11076 22332
rect 11132 22330 11156 22332
rect 11212 22330 11236 22332
rect 10972 22278 10982 22330
rect 11226 22278 11236 22330
rect 10972 22276 10996 22278
rect 11052 22276 11076 22278
rect 11132 22276 11156 22278
rect 11212 22276 11236 22278
rect 10916 22267 11292 22276
rect 11992 22094 12020 22578
rect 11992 22066 12112 22094
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11164 21690 11192 21898
rect 11656 21788 12032 21797
rect 11712 21786 11736 21788
rect 11792 21786 11816 21788
rect 11872 21786 11896 21788
rect 11952 21786 11976 21788
rect 11712 21734 11722 21786
rect 11966 21734 11976 21786
rect 11712 21732 11736 21734
rect 11792 21732 11816 21734
rect 11872 21732 11896 21734
rect 11952 21732 11976 21734
rect 11656 21723 12032 21732
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 10916 21244 11292 21253
rect 10972 21242 10996 21244
rect 11052 21242 11076 21244
rect 11132 21242 11156 21244
rect 11212 21242 11236 21244
rect 10972 21190 10982 21242
rect 11226 21190 11236 21242
rect 10972 21188 10996 21190
rect 11052 21188 11076 21190
rect 11132 21188 11156 21190
rect 11212 21188 11236 21190
rect 10916 21179 11292 21188
rect 11656 20700 12032 20709
rect 11712 20698 11736 20700
rect 11792 20698 11816 20700
rect 11872 20698 11896 20700
rect 11952 20698 11976 20700
rect 11712 20646 11722 20698
rect 11966 20646 11976 20698
rect 11712 20644 11736 20646
rect 11792 20644 11816 20646
rect 11872 20644 11896 20646
rect 11952 20644 11976 20646
rect 11656 20635 12032 20644
rect 10916 20156 11292 20165
rect 10972 20154 10996 20156
rect 11052 20154 11076 20156
rect 11132 20154 11156 20156
rect 11212 20154 11236 20156
rect 10972 20102 10982 20154
rect 11226 20102 11236 20154
rect 10972 20100 10996 20102
rect 11052 20100 11076 20102
rect 11132 20100 11156 20102
rect 11212 20100 11236 20102
rect 10916 20091 11292 20100
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10980 19446 11008 19790
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11532 19514 11560 19722
rect 11656 19612 12032 19621
rect 11712 19610 11736 19612
rect 11792 19610 11816 19612
rect 11872 19610 11896 19612
rect 11952 19610 11976 19612
rect 11712 19558 11722 19610
rect 11966 19558 11976 19610
rect 11712 19556 11736 19558
rect 11792 19556 11816 19558
rect 11872 19556 11896 19558
rect 11952 19556 11976 19558
rect 11656 19547 12032 19556
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10704 18902 10732 19246
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 10916 19068 11292 19077
rect 10972 19066 10996 19068
rect 11052 19066 11076 19068
rect 11132 19066 11156 19068
rect 11212 19066 11236 19068
rect 10972 19014 10982 19066
rect 11226 19014 11236 19066
rect 10972 19012 10996 19014
rect 11052 19012 11076 19014
rect 11132 19012 11156 19014
rect 11212 19012 11236 19014
rect 10916 19003 11292 19012
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10428 17870 10548 17898
rect 10600 17876 10652 17882
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10244 14906 10272 17206
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10336 16590 10364 16934
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10336 15706 10364 16050
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10336 15162 10364 15642
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10244 14878 10364 14906
rect 10336 14362 10364 14878
rect 10244 14334 10364 14362
rect 10244 12850 10272 14334
rect 10428 13802 10456 17870
rect 10600 17818 10652 17824
rect 10612 17678 10640 17818
rect 10796 17746 10824 18906
rect 10916 17980 11292 17989
rect 10972 17978 10996 17980
rect 11052 17978 11076 17980
rect 11132 17978 11156 17980
rect 11212 17978 11236 17980
rect 10972 17926 10982 17978
rect 11226 17926 11236 17978
rect 10972 17924 10996 17926
rect 11052 17924 11076 17926
rect 11132 17924 11156 17926
rect 11212 17924 11236 17926
rect 10916 17915 11292 17924
rect 11440 17814 11468 19178
rect 11900 18766 11928 19314
rect 12084 18970 12112 22066
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12268 20534 12296 21490
rect 12360 21486 12388 25298
rect 12452 23662 12480 26318
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 23254 12480 23598
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12452 22030 12480 23190
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 12176 19378 12204 19654
rect 12268 19514 12296 20470
rect 12544 19938 12572 26998
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12728 26382 12756 26726
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 13004 25498 13032 26930
rect 13360 26784 13412 26790
rect 13360 26726 13412 26732
rect 13372 25974 13400 26726
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 12808 23792 12860 23798
rect 12808 23734 12860 23740
rect 12820 23594 12848 23734
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 13188 23118 13216 24006
rect 13176 23112 13228 23118
rect 12898 23080 12954 23089
rect 13176 23054 13228 23060
rect 12898 23015 12900 23024
rect 12952 23015 12954 23024
rect 12900 22986 12952 22992
rect 12912 22710 12940 22986
rect 13372 22778 13400 24142
rect 13464 23866 13492 25094
rect 13556 24818 13584 26930
rect 13820 26920 13872 26926
rect 13820 26862 13872 26868
rect 13832 26246 13860 26862
rect 14476 26858 14504 27406
rect 15656 27228 16032 27237
rect 15712 27226 15736 27228
rect 15792 27226 15816 27228
rect 15872 27226 15896 27228
rect 15952 27226 15976 27228
rect 15712 27174 15722 27226
rect 15966 27174 15976 27226
rect 15712 27172 15736 27174
rect 15792 27172 15816 27174
rect 15872 27172 15896 27174
rect 15952 27172 15976 27174
rect 15656 27163 16032 27172
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 14464 26852 14516 26858
rect 14464 26794 14516 26800
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13832 25294 13860 26182
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 12900 22704 12952 22710
rect 12900 22646 12952 22652
rect 13464 22642 13492 23802
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13556 22574 13584 24074
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13740 22778 13768 22918
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 12636 22234 12664 22510
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 12636 21690 12664 22170
rect 12728 22166 12756 22374
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12452 19910 12572 19938
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 11656 18524 12032 18533
rect 11712 18522 11736 18524
rect 11792 18522 11816 18524
rect 11872 18522 11896 18524
rect 11952 18522 11976 18524
rect 11712 18470 11722 18522
rect 11966 18470 11976 18522
rect 11712 18468 11736 18470
rect 11792 18468 11816 18470
rect 11872 18468 11896 18470
rect 11952 18468 11976 18470
rect 11656 18459 12032 18468
rect 12084 18222 12112 18702
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 12268 17746 12296 19450
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10520 16250 10548 17138
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10508 15496 10560 15502
rect 10506 15464 10508 15473
rect 10560 15464 10562 15473
rect 10506 15399 10562 15408
rect 10612 15026 10640 17614
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10704 16794 10732 17546
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 10916 16892 11292 16901
rect 10972 16890 10996 16892
rect 11052 16890 11076 16892
rect 11132 16890 11156 16892
rect 11212 16890 11236 16892
rect 10972 16838 10982 16890
rect 11226 16838 11236 16890
rect 10972 16836 10996 16838
rect 11052 16836 11076 16838
rect 11132 16836 11156 16838
rect 11212 16836 11236 16838
rect 10916 16827 11292 16836
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10704 16250 10732 16730
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10980 16046 11008 16662
rect 11348 16590 11376 17478
rect 11656 17436 12032 17445
rect 11712 17434 11736 17436
rect 11792 17434 11816 17436
rect 11872 17434 11896 17436
rect 11952 17434 11976 17436
rect 11712 17382 11722 17434
rect 11966 17382 11976 17434
rect 11712 17380 11736 17382
rect 11792 17380 11816 17382
rect 11872 17380 11896 17382
rect 11952 17380 11976 17382
rect 11656 17371 12032 17380
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11532 16590 11560 16934
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11440 16114 11468 16390
rect 11656 16348 12032 16357
rect 11712 16346 11736 16348
rect 11792 16346 11816 16348
rect 11872 16346 11896 16348
rect 11952 16346 11976 16348
rect 11712 16294 11722 16346
rect 11966 16294 11976 16346
rect 11712 16292 11736 16294
rect 11792 16292 11816 16294
rect 11872 16292 11896 16294
rect 11952 16292 11976 16294
rect 11656 16283 12032 16292
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 10876 16040 10928 16046
rect 10874 16008 10876 16017
rect 10968 16040 11020 16046
rect 10928 16008 10930 16017
rect 10968 15982 11020 15988
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 10874 15943 10930 15952
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 10916 15804 11292 15813
rect 10972 15802 10996 15804
rect 11052 15802 11076 15804
rect 11132 15802 11156 15804
rect 11212 15802 11236 15804
rect 10972 15750 10982 15802
rect 11226 15750 11236 15802
rect 10972 15748 10996 15750
rect 11052 15748 11076 15750
rect 11132 15748 11156 15750
rect 11212 15748 11236 15750
rect 10916 15739 11292 15748
rect 11348 15502 11376 15914
rect 11716 15570 11744 15982
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 10888 15162 10916 15438
rect 12268 15434 12296 16458
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11656 15260 12032 15269
rect 11712 15258 11736 15260
rect 11792 15258 11816 15260
rect 11872 15258 11896 15260
rect 11952 15258 11976 15260
rect 11712 15206 11722 15258
rect 11966 15206 11976 15258
rect 11712 15204 11736 15206
rect 11792 15204 11816 15206
rect 11872 15204 11896 15206
rect 11952 15204 11976 15206
rect 11058 15192 11114 15201
rect 11656 15195 12032 15204
rect 10876 15156 10928 15162
rect 11058 15127 11060 15136
rect 10876 15098 10928 15104
rect 11112 15127 11114 15136
rect 11428 15156 11480 15162
rect 11060 15098 11112 15104
rect 11428 15098 11480 15104
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10916 14716 11292 14725
rect 10972 14714 10996 14716
rect 11052 14714 11076 14716
rect 11132 14714 11156 14716
rect 11212 14714 11236 14716
rect 10972 14662 10982 14714
rect 11226 14662 11236 14714
rect 10972 14660 10996 14662
rect 11052 14660 11076 14662
rect 11132 14660 11156 14662
rect 11212 14660 11236 14662
rect 10916 14651 11292 14660
rect 11440 13938 11468 15098
rect 12084 14550 12112 15302
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 11656 14172 12032 14181
rect 11712 14170 11736 14172
rect 11792 14170 11816 14172
rect 11872 14170 11896 14172
rect 11952 14170 11976 14172
rect 11712 14118 11722 14170
rect 11966 14118 11976 14170
rect 11712 14116 11736 14118
rect 11792 14116 11816 14118
rect 11872 14116 11896 14118
rect 11952 14116 11976 14118
rect 11656 14107 12032 14116
rect 12084 13938 12112 14486
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10232 12640 10284 12646
rect 10284 12600 10364 12628
rect 10232 12582 10284 12588
rect 10336 11762 10364 12600
rect 10520 12306 10548 13126
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11830 10548 12038
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10046 10775 10048 10784
rect 10100 10775 10102 10784
rect 10140 10804 10192 10810
rect 10048 10746 10100 10752
rect 10140 10746 10192 10752
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10152 9518 10180 9658
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10152 7478 10180 9454
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6322 9812 6598
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8864 5902 8984 5930
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 7656 5468 8032 5477
rect 7712 5466 7736 5468
rect 7792 5466 7816 5468
rect 7872 5466 7896 5468
rect 7952 5466 7976 5468
rect 7712 5414 7722 5466
rect 7966 5414 7976 5466
rect 7712 5412 7736 5414
rect 7792 5412 7816 5414
rect 7872 5412 7896 5414
rect 7952 5412 7976 5414
rect 7656 5403 8032 5412
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7944 4690 7972 5238
rect 8128 5234 8156 5510
rect 8220 5370 8248 5850
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7656 4380 8032 4389
rect 7712 4378 7736 4380
rect 7792 4378 7816 4380
rect 7872 4378 7896 4380
rect 7952 4378 7976 4380
rect 7712 4326 7722 4378
rect 7966 4326 7976 4378
rect 7712 4324 7736 4326
rect 7792 4324 7816 4326
rect 7872 4324 7896 4326
rect 7952 4324 7976 4326
rect 7656 4315 8032 4324
rect 8220 3738 8248 5034
rect 8312 4554 8340 5102
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8312 4282 8340 4490
rect 8404 4486 8432 5646
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8404 4146 8432 4422
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 7656 3292 8032 3301
rect 7712 3290 7736 3292
rect 7792 3290 7816 3292
rect 7872 3290 7896 3292
rect 7952 3290 7976 3292
rect 7712 3238 7722 3290
rect 7966 3238 7976 3290
rect 7712 3236 7736 3238
rect 7792 3236 7816 3238
rect 7872 3236 7896 3238
rect 7952 3236 7976 3238
rect 7656 3227 8032 3236
rect 8220 3194 8248 3674
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8404 3058 8432 4082
rect 8864 4078 8892 5902
rect 9048 5370 9076 6190
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8864 3466 8892 4014
rect 8956 3534 8984 4966
rect 9232 4826 9260 6258
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5166 9444 5510
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 4282 9168 4558
rect 9416 4554 9444 5102
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 3126 9168 3334
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 9232 3058 9260 3538
rect 9324 3534 9352 4422
rect 9508 4146 9536 6258
rect 9876 5914 9904 6734
rect 10244 6458 10272 10542
rect 10428 10266 10456 10610
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10336 9450 10364 10202
rect 10428 9722 10456 10202
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10324 9444 10376 9450
rect 10324 9386 10376 9392
rect 10520 8634 10548 10610
rect 10612 9738 10640 13330
rect 10704 13326 10732 13874
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 10916 13628 11292 13637
rect 10972 13626 10996 13628
rect 11052 13626 11076 13628
rect 11132 13626 11156 13628
rect 11212 13626 11236 13628
rect 10972 13574 10982 13626
rect 11226 13574 11236 13626
rect 10972 13572 10996 13574
rect 11052 13572 11076 13574
rect 11132 13572 11156 13574
rect 11212 13572 11236 13574
rect 10916 13563 11292 13572
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12986 10732 13262
rect 11348 13258 11376 13670
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 11072 12850 11100 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10916 12540 11292 12549
rect 10972 12538 10996 12540
rect 11052 12538 11076 12540
rect 11132 12538 11156 12540
rect 11212 12538 11236 12540
rect 10972 12486 10982 12538
rect 11226 12486 11236 12538
rect 10972 12484 10996 12486
rect 11052 12484 11076 12486
rect 11132 12484 11156 12486
rect 11212 12484 11236 12486
rect 10916 12475 11292 12484
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10704 11830 10732 12106
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 10916 11452 11292 11461
rect 10972 11450 10996 11452
rect 11052 11450 11076 11452
rect 11132 11450 11156 11452
rect 11212 11450 11236 11452
rect 10972 11398 10982 11450
rect 11226 11398 11236 11450
rect 10972 11396 10996 11398
rect 11052 11396 11076 11398
rect 11132 11396 11156 11398
rect 11212 11396 11236 11398
rect 10916 11387 11292 11396
rect 10916 10364 11292 10373
rect 10972 10362 10996 10364
rect 11052 10362 11076 10364
rect 11132 10362 11156 10364
rect 11212 10362 11236 10364
rect 10972 10310 10982 10362
rect 11226 10310 11236 10362
rect 10972 10308 10996 10310
rect 11052 10308 11076 10310
rect 11132 10308 11156 10310
rect 11212 10308 11236 10310
rect 10916 10299 11292 10308
rect 10612 9710 10732 9738
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 8906 10640 9522
rect 10704 9450 10732 9710
rect 11348 9450 11376 11698
rect 11440 10810 11468 13874
rect 11808 13530 11836 13874
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11532 12986 11560 13466
rect 11656 13084 12032 13093
rect 11712 13082 11736 13084
rect 11792 13082 11816 13084
rect 11872 13082 11896 13084
rect 11952 13082 11976 13084
rect 11712 13030 11722 13082
rect 11966 13030 11976 13082
rect 11712 13028 11736 13030
rect 11792 13028 11816 13030
rect 11872 13028 11896 13030
rect 11952 13028 11976 13030
rect 11656 13019 12032 13028
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10248 11560 12718
rect 12084 12434 12112 13874
rect 12176 12986 12204 13874
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12084 12406 12204 12434
rect 11656 11996 12032 12005
rect 11712 11994 11736 11996
rect 11792 11994 11816 11996
rect 11872 11994 11896 11996
rect 11952 11994 11976 11996
rect 11712 11942 11722 11994
rect 11966 11942 11976 11994
rect 11712 11940 11736 11942
rect 11792 11940 11816 11942
rect 11872 11940 11896 11942
rect 11952 11940 11976 11942
rect 11656 11931 12032 11940
rect 12176 11082 12204 12406
rect 12268 11898 12296 13806
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11656 10908 12032 10917
rect 11712 10906 11736 10908
rect 11792 10906 11816 10908
rect 11872 10906 11896 10908
rect 11952 10906 11976 10908
rect 11712 10854 11722 10906
rect 11966 10854 11976 10906
rect 11712 10852 11736 10854
rect 11792 10852 11816 10854
rect 11872 10852 11896 10854
rect 11952 10852 11976 10854
rect 11656 10843 12032 10852
rect 11440 10220 11560 10248
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10612 8537 10640 8842
rect 10598 8528 10654 8537
rect 10598 8463 10654 8472
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10336 7206 10364 7278
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10244 5710 10272 6394
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9784 4622 9812 5170
rect 10336 4690 10364 7142
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9508 3738 9536 4082
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9784 3194 9812 4558
rect 10612 4486 10640 7346
rect 10704 5778 10732 9386
rect 10916 9276 11292 9285
rect 10972 9274 10996 9276
rect 11052 9274 11076 9276
rect 11132 9274 11156 9276
rect 11212 9274 11236 9276
rect 10972 9222 10982 9274
rect 11226 9222 11236 9274
rect 10972 9220 10996 9222
rect 11052 9220 11076 9222
rect 11132 9220 11156 9222
rect 11212 9220 11236 9222
rect 10916 9211 11292 9220
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8498 10824 8774
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10916 8188 11292 8197
rect 10972 8186 10996 8188
rect 11052 8186 11076 8188
rect 11132 8186 11156 8188
rect 11212 8186 11236 8188
rect 10972 8134 10982 8186
rect 11226 8134 11236 8186
rect 10972 8132 10996 8134
rect 11052 8132 11076 8134
rect 11132 8132 11156 8134
rect 11212 8132 11236 8134
rect 10916 8123 11292 8132
rect 11348 7886 11376 9386
rect 11440 9382 11468 10220
rect 12084 9994 12112 10950
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 11656 9820 12032 9829
rect 11712 9818 11736 9820
rect 11792 9818 11816 9820
rect 11872 9818 11896 9820
rect 11952 9818 11976 9820
rect 11712 9766 11722 9818
rect 11966 9766 11976 9818
rect 11712 9764 11736 9766
rect 11792 9764 11816 9766
rect 11872 9764 11896 9766
rect 11952 9764 11976 9766
rect 11656 9755 12032 9764
rect 12176 9654 12204 11018
rect 12452 9926 12480 19910
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 19378 12572 19790
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12820 17542 12848 20538
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 19446 13124 20198
rect 13280 20058 13308 20402
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 13372 19854 13400 20198
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12636 16250 12664 17070
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12636 15910 12664 16186
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13326 12572 13670
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12728 11218 12756 14418
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10266 12756 10950
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11440 8838 11468 9318
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11656 8732 12032 8741
rect 11712 8730 11736 8732
rect 11792 8730 11816 8732
rect 11872 8730 11896 8732
rect 11952 8730 11976 8732
rect 11712 8678 11722 8730
rect 11966 8678 11976 8730
rect 11712 8676 11736 8678
rect 11792 8676 11816 8678
rect 11872 8676 11896 8678
rect 11952 8676 11976 8678
rect 11656 8667 12032 8676
rect 12176 8498 12204 9590
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12452 8838 12480 9114
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12636 8498 12664 8910
rect 12820 8906 12848 17478
rect 13004 17338 13032 18634
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12900 17128 12952 17134
rect 12898 17096 12900 17105
rect 12952 17096 12954 17105
rect 12898 17031 12954 17040
rect 13188 16590 13216 17614
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16794 13308 17138
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13188 16096 13216 16526
rect 13096 16068 13216 16096
rect 13096 15910 13124 16068
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12918 13124 13126
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13280 12442 13308 13262
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13372 12102 13400 19654
rect 13464 14482 13492 20334
rect 13556 19514 13584 20402
rect 13648 19786 13676 22578
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13740 20466 13768 22374
rect 13924 22166 13952 26726
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14108 25820 14136 26318
rect 14280 25832 14332 25838
rect 14108 25792 14280 25820
rect 14108 23118 14136 25792
rect 14280 25774 14332 25780
rect 14476 25770 14504 26794
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14660 25974 14688 26726
rect 14752 26314 14780 26726
rect 14740 26308 14792 26314
rect 14740 26250 14792 26256
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14464 25764 14516 25770
rect 14464 25706 14516 25712
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 13912 22160 13964 22166
rect 13912 22102 13964 22108
rect 14108 21554 14136 23054
rect 14292 22506 14320 23462
rect 14844 23322 14872 26930
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16488 26784 16540 26790
rect 16488 26726 16540 26732
rect 14916 26684 15292 26693
rect 14972 26682 14996 26684
rect 15052 26682 15076 26684
rect 15132 26682 15156 26684
rect 15212 26682 15236 26684
rect 14972 26630 14982 26682
rect 15226 26630 15236 26682
rect 14972 26628 14996 26630
rect 15052 26628 15076 26630
rect 15132 26628 15156 26630
rect 15212 26628 15236 26630
rect 14916 26619 15292 26628
rect 16500 26314 16528 26726
rect 15568 26308 15620 26314
rect 15568 26250 15620 26256
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 15580 26042 15608 26250
rect 16120 26240 16172 26246
rect 16120 26182 16172 26188
rect 15656 26140 16032 26149
rect 15712 26138 15736 26140
rect 15792 26138 15816 26140
rect 15872 26138 15896 26140
rect 15952 26138 15976 26140
rect 15712 26086 15722 26138
rect 15966 26086 15976 26138
rect 15712 26084 15736 26086
rect 15792 26084 15816 26086
rect 15872 26084 15896 26086
rect 15952 26084 15976 26086
rect 15656 26075 16032 26084
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 14916 25596 15292 25605
rect 14972 25594 14996 25596
rect 15052 25594 15076 25596
rect 15132 25594 15156 25596
rect 15212 25594 15236 25596
rect 14972 25542 14982 25594
rect 15226 25542 15236 25594
rect 14972 25540 14996 25542
rect 15052 25540 15076 25542
rect 15132 25540 15156 25542
rect 15212 25540 15236 25542
rect 14916 25531 15292 25540
rect 15396 25498 15424 25910
rect 16132 25906 16160 26182
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15656 25052 16032 25061
rect 15712 25050 15736 25052
rect 15792 25050 15816 25052
rect 15872 25050 15896 25052
rect 15952 25050 15976 25052
rect 15712 24998 15722 25050
rect 15966 24998 15976 25050
rect 15712 24996 15736 24998
rect 15792 24996 15816 24998
rect 15872 24996 15896 24998
rect 15952 24996 15976 24998
rect 15656 24987 16032 24996
rect 15568 24948 15620 24954
rect 15568 24890 15620 24896
rect 15580 24818 15608 24890
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 14916 24508 15292 24517
rect 14972 24506 14996 24508
rect 15052 24506 15076 24508
rect 15132 24506 15156 24508
rect 15212 24506 15236 24508
rect 14972 24454 14982 24506
rect 15226 24454 15236 24506
rect 14972 24452 14996 24454
rect 15052 24452 15076 24454
rect 15132 24452 15156 24454
rect 15212 24452 15236 24454
rect 14916 24443 15292 24452
rect 15580 23662 15608 24754
rect 15656 23964 16032 23973
rect 15712 23962 15736 23964
rect 15792 23962 15816 23964
rect 15872 23962 15896 23964
rect 15952 23962 15976 23964
rect 15712 23910 15722 23962
rect 15966 23910 15976 23962
rect 15712 23908 15736 23910
rect 15792 23908 15816 23910
rect 15872 23908 15896 23910
rect 15952 23908 15976 23910
rect 15656 23899 16032 23908
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 14916 23420 15292 23429
rect 14972 23418 14996 23420
rect 15052 23418 15076 23420
rect 15132 23418 15156 23420
rect 15212 23418 15236 23420
rect 14972 23366 14982 23418
rect 15226 23366 15236 23418
rect 14972 23364 14996 23366
rect 15052 23364 15076 23366
rect 15132 23364 15156 23366
rect 15212 23364 15236 23366
rect 14916 23355 15292 23364
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 16132 23118 16160 25842
rect 16592 25770 16620 26862
rect 17236 26790 17264 26930
rect 17408 26920 17460 26926
rect 17328 26868 17408 26874
rect 17328 26862 17460 26868
rect 17328 26846 17448 26862
rect 17500 26852 17552 26858
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 26042 16712 26522
rect 17328 26042 17356 26846
rect 17500 26794 17552 26800
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 17316 26036 17368 26042
rect 17316 25978 17368 25984
rect 16580 25764 16632 25770
rect 16580 25706 16632 25712
rect 16304 25696 16356 25702
rect 16304 25638 16356 25644
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16316 25226 16344 25638
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14384 22778 14412 22986
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15488 22778 15516 22918
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13740 17202 13768 19926
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13636 16584 13688 16590
rect 13634 16552 13636 16561
rect 13688 16552 13690 16561
rect 13544 16516 13596 16522
rect 13634 16487 13690 16496
rect 13544 16458 13596 16464
rect 13556 16114 13584 16458
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13556 15706 13584 16050
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13450 14376 13506 14385
rect 13450 14311 13506 14320
rect 13464 13376 13492 14311
rect 13544 13796 13596 13802
rect 13648 13784 13676 16487
rect 13740 14618 13768 17138
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16794 13860 17070
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13596 13756 13676 13784
rect 13544 13738 13596 13744
rect 13464 13348 13584 13376
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 12912 11014 12940 12038
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10606 12940 10950
rect 13188 10810 13216 11018
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12820 8566 12848 8842
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11440 8090 11468 8366
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11428 7948 11480 7954
rect 11612 7948 11664 7954
rect 11428 7890 11480 7896
rect 11532 7908 11612 7936
rect 11336 7880 11388 7886
rect 11242 7848 11298 7857
rect 11336 7822 11388 7828
rect 11242 7783 11298 7792
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7546 10824 7686
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 7290 11008 7346
rect 10796 7262 11008 7290
rect 11256 7274 11284 7783
rect 11244 7268 11296 7274
rect 10796 7002 10824 7262
rect 11244 7210 11296 7216
rect 10916 7100 11292 7109
rect 10972 7098 10996 7100
rect 11052 7098 11076 7100
rect 11132 7098 11156 7100
rect 11212 7098 11236 7100
rect 10972 7046 10982 7098
rect 11226 7046 11236 7098
rect 10972 7044 10996 7046
rect 11052 7044 11076 7046
rect 11132 7044 11156 7046
rect 11212 7044 11236 7046
rect 10916 7035 11292 7044
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10916 6012 11292 6021
rect 10972 6010 10996 6012
rect 11052 6010 11076 6012
rect 11132 6010 11156 6012
rect 11212 6010 11236 6012
rect 10972 5958 10982 6010
rect 11226 5958 11236 6010
rect 10972 5956 10996 5958
rect 11052 5956 11076 5958
rect 11132 5956 11156 5958
rect 11212 5956 11236 5958
rect 10916 5947 11292 5956
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10916 4924 11292 4933
rect 10972 4922 10996 4924
rect 11052 4922 11076 4924
rect 11132 4922 11156 4924
rect 11212 4922 11236 4924
rect 10972 4870 10982 4922
rect 11226 4870 11236 4922
rect 10972 4868 10996 4870
rect 11052 4868 11076 4870
rect 11132 4868 11156 4870
rect 11212 4868 11236 4870
rect 10916 4859 11292 4868
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10244 3942 10272 4422
rect 10704 4282 10732 4626
rect 10796 4554 11008 4570
rect 10784 4548 11020 4554
rect 10836 4542 10968 4548
rect 10784 4490 10836 4496
rect 10968 4490 11020 4496
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10612 3942 10640 4082
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10704 3670 10732 4218
rect 11164 4146 11192 4694
rect 11348 4486 11376 7822
rect 11440 7002 11468 7890
rect 11532 7342 11560 7908
rect 11612 7890 11664 7896
rect 11716 7886 11744 8230
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11656 7644 12032 7653
rect 11712 7642 11736 7644
rect 11792 7642 11816 7644
rect 11872 7642 11896 7644
rect 11952 7642 11976 7644
rect 11712 7590 11722 7642
rect 11966 7590 11976 7642
rect 11712 7588 11736 7590
rect 11792 7588 11816 7590
rect 11872 7588 11896 7590
rect 11952 7588 11976 7590
rect 11656 7579 12032 7588
rect 12084 7478 12112 8026
rect 12636 7546 12664 8434
rect 12716 8424 12768 8430
rect 12912 8378 12940 10542
rect 12768 8372 12940 8378
rect 12716 8366 12940 8372
rect 12728 8350 12940 8366
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11532 6254 11560 7278
rect 11656 6556 12032 6565
rect 11712 6554 11736 6556
rect 11792 6554 11816 6556
rect 11872 6554 11896 6556
rect 11952 6554 11976 6556
rect 11712 6502 11722 6554
rect 11966 6502 11976 6554
rect 11712 6500 11736 6502
rect 11792 6500 11816 6502
rect 11872 6500 11896 6502
rect 11952 6500 11976 6502
rect 11656 6491 12032 6500
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11808 5914 11836 6258
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 12728 5846 12756 8350
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 13004 5710 13032 6054
rect 13188 5914 13216 10610
rect 13464 10062 13492 10746
rect 13556 10062 13584 13348
rect 13648 10112 13676 13756
rect 13740 10674 13768 14418
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13394 13860 13670
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13924 11506 13952 20198
rect 14016 19854 14044 20402
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14016 19378 14044 19790
rect 14108 19446 14136 21490
rect 14476 21146 14504 21490
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14108 18834 14136 19382
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14004 17740 14056 17746
rect 14200 17728 14228 19858
rect 14292 19718 14320 20266
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14292 19514 14320 19654
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14056 17700 14228 17728
rect 14004 17682 14056 17688
rect 14016 16046 14044 17682
rect 14292 16538 14320 19110
rect 14384 18766 14412 20402
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14660 19514 14688 19722
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14384 17202 14412 17614
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14384 16590 14412 17138
rect 14108 16510 14320 16538
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14004 15088 14056 15094
rect 14002 15056 14004 15065
rect 14056 15056 14058 15065
rect 14002 14991 14058 15000
rect 14108 12850 14136 16510
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16182 14320 16390
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14200 15706 14228 16050
rect 14384 16046 14412 16526
rect 14568 16250 14596 17138
rect 14752 16454 14780 18158
rect 14844 18154 14872 22442
rect 14916 22332 15292 22341
rect 14972 22330 14996 22332
rect 15052 22330 15076 22332
rect 15132 22330 15156 22332
rect 15212 22330 15236 22332
rect 14972 22278 14982 22330
rect 15226 22278 15236 22330
rect 14972 22276 14996 22278
rect 15052 22276 15076 22278
rect 15132 22276 15156 22278
rect 15212 22276 15236 22278
rect 14916 22267 15292 22276
rect 15488 22098 15516 22714
rect 15580 22234 15608 23054
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 15656 22876 16032 22885
rect 15712 22874 15736 22876
rect 15792 22874 15816 22876
rect 15872 22874 15896 22876
rect 15952 22874 15976 22876
rect 15712 22822 15722 22874
rect 15966 22822 15976 22874
rect 15712 22820 15736 22822
rect 15792 22820 15816 22822
rect 15872 22820 15896 22822
rect 15952 22820 15976 22822
rect 15656 22811 16032 22820
rect 16132 22642 16160 22918
rect 16224 22710 16252 25094
rect 16316 23118 16344 25162
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 16212 22704 16264 22710
rect 16212 22646 16264 22652
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15476 21956 15528 21962
rect 15476 21898 15528 21904
rect 14916 21244 15292 21253
rect 14972 21242 14996 21244
rect 15052 21242 15076 21244
rect 15132 21242 15156 21244
rect 15212 21242 15236 21244
rect 14972 21190 14982 21242
rect 15226 21190 15236 21242
rect 14972 21188 14996 21190
rect 15052 21188 15076 21190
rect 15132 21188 15156 21190
rect 15212 21188 15236 21190
rect 14916 21179 15292 21188
rect 15396 20602 15424 21898
rect 15488 21690 15516 21898
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15580 21350 15608 21966
rect 15656 21788 16032 21797
rect 15712 21786 15736 21788
rect 15792 21786 15816 21788
rect 15872 21786 15896 21788
rect 15952 21786 15976 21788
rect 15712 21734 15722 21786
rect 15966 21734 15976 21786
rect 15712 21732 15736 21734
rect 15792 21732 15816 21734
rect 15872 21732 15896 21734
rect 15952 21732 15976 21734
rect 15656 21723 16032 21732
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15580 20890 15608 21286
rect 15672 20942 15700 21286
rect 15488 20862 15608 20890
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15488 20369 15516 20862
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15474 20360 15530 20369
rect 15474 20295 15530 20304
rect 14916 20156 15292 20165
rect 14972 20154 14996 20156
rect 15052 20154 15076 20156
rect 15132 20154 15156 20156
rect 15212 20154 15236 20156
rect 14972 20102 14982 20154
rect 15226 20102 15236 20154
rect 14972 20100 14996 20102
rect 15052 20100 15076 20102
rect 15132 20100 15156 20102
rect 15212 20100 15236 20102
rect 14916 20091 15292 20100
rect 14916 19068 15292 19077
rect 14972 19066 14996 19068
rect 15052 19066 15076 19068
rect 15132 19066 15156 19068
rect 15212 19066 15236 19068
rect 14972 19014 14982 19066
rect 15226 19014 15236 19066
rect 14972 19012 14996 19014
rect 15052 19012 15076 19014
rect 15132 19012 15156 19014
rect 15212 19012 15236 19014
rect 14916 19003 15292 19012
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15120 18426 15148 18634
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14844 16658 14872 18090
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 14916 17980 15292 17989
rect 14972 17978 14996 17980
rect 15052 17978 15076 17980
rect 15132 17978 15156 17980
rect 15212 17978 15236 17980
rect 14972 17926 14982 17978
rect 15226 17926 15236 17978
rect 14972 17924 14996 17926
rect 15052 17924 15076 17926
rect 15132 17924 15156 17926
rect 15212 17924 15236 17926
rect 14916 17915 15292 17924
rect 14916 16892 15292 16901
rect 14972 16890 14996 16892
rect 15052 16890 15076 16892
rect 15132 16890 15156 16892
rect 15212 16890 15236 16892
rect 14972 16838 14982 16890
rect 15226 16838 15236 16890
rect 14972 16836 14996 16838
rect 15052 16836 15076 16838
rect 15132 16836 15156 16838
rect 15212 16836 15236 16838
rect 14916 16827 15292 16836
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14844 16130 14872 16594
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14568 16102 14872 16130
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14200 13258 14228 14010
rect 14292 14006 14320 14214
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14384 13734 14412 15982
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14476 12986 14504 13874
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14016 12170 14044 12582
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 14016 11762 14044 12106
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14464 11552 14516 11558
rect 13924 11478 14044 11506
rect 14464 11494 14516 11500
rect 14016 10674 14044 11478
rect 14476 10674 14504 11494
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 14568 10146 14596 16102
rect 14936 15994 14964 16390
rect 14752 15966 14964 15994
rect 14752 15366 14780 15966
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14844 15502 14872 15846
rect 14916 15804 15292 15813
rect 14972 15802 14996 15804
rect 15052 15802 15076 15804
rect 15132 15802 15156 15804
rect 15212 15802 15236 15804
rect 14972 15750 14982 15802
rect 15226 15750 15236 15802
rect 14972 15748 14996 15750
rect 15052 15748 15076 15750
rect 15132 15748 15156 15750
rect 15212 15748 15236 15750
rect 14916 15739 15292 15748
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14752 14260 14780 15302
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14844 14521 14872 14758
rect 14916 14716 15292 14725
rect 14972 14714 14996 14716
rect 15052 14714 15076 14716
rect 15132 14714 15156 14716
rect 15212 14714 15236 14716
rect 14972 14662 14982 14714
rect 15226 14662 15236 14714
rect 14972 14660 14996 14662
rect 15052 14660 15076 14662
rect 15132 14660 15156 14662
rect 15212 14660 15236 14662
rect 14916 14651 15292 14660
rect 14830 14512 14886 14521
rect 15396 14498 15424 18022
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15488 15434 15516 16934
rect 15580 16697 15608 20742
rect 15656 20700 16032 20709
rect 15712 20698 15736 20700
rect 15792 20698 15816 20700
rect 15872 20698 15896 20700
rect 15952 20698 15976 20700
rect 15712 20646 15722 20698
rect 15966 20646 15976 20698
rect 15712 20644 15736 20646
rect 15792 20644 15816 20646
rect 15872 20644 15896 20646
rect 15952 20644 15976 20646
rect 15656 20635 16032 20644
rect 15656 19612 16032 19621
rect 15712 19610 15736 19612
rect 15792 19610 15816 19612
rect 15872 19610 15896 19612
rect 15952 19610 15976 19612
rect 15712 19558 15722 19610
rect 15966 19558 15976 19610
rect 15712 19556 15736 19558
rect 15792 19556 15816 19558
rect 15872 19556 15896 19558
rect 15952 19556 15976 19558
rect 15656 19547 16032 19556
rect 15656 18524 16032 18533
rect 15712 18522 15736 18524
rect 15792 18522 15816 18524
rect 15872 18522 15896 18524
rect 15952 18522 15976 18524
rect 15712 18470 15722 18522
rect 15966 18470 15976 18522
rect 15712 18468 15736 18470
rect 15792 18468 15816 18470
rect 15872 18468 15896 18470
rect 15952 18468 15976 18470
rect 15656 18459 16032 18468
rect 16132 18154 16160 22578
rect 16224 22094 16252 22646
rect 16224 22066 16344 22094
rect 16316 21554 16344 22066
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15656 17436 16032 17445
rect 15712 17434 15736 17436
rect 15792 17434 15816 17436
rect 15872 17434 15896 17436
rect 15952 17434 15976 17436
rect 15712 17382 15722 17434
rect 15966 17382 15976 17434
rect 15712 17380 15736 17382
rect 15792 17380 15816 17382
rect 15872 17380 15896 17382
rect 15952 17380 15976 17382
rect 15656 17371 16032 17380
rect 16132 17202 16160 17478
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15566 16688 15622 16697
rect 15566 16623 15622 16632
rect 16040 16590 16068 17138
rect 16028 16584 16080 16590
rect 16080 16532 16160 16538
rect 16028 16526 16160 16532
rect 15568 16516 15620 16522
rect 16040 16510 16160 16526
rect 15568 16458 15620 16464
rect 15580 16250 15608 16458
rect 15656 16348 16032 16357
rect 15712 16346 15736 16348
rect 15792 16346 15816 16348
rect 15872 16346 15896 16348
rect 15952 16346 15976 16348
rect 15712 16294 15722 16346
rect 15966 16294 15976 16346
rect 15712 16292 15736 16294
rect 15792 16292 15816 16294
rect 15872 16292 15896 16294
rect 15952 16292 15976 16294
rect 15656 16283 16032 16292
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15580 15570 15608 16050
rect 16132 15978 16160 16510
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15396 14470 15516 14498
rect 14830 14447 14886 14456
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 14832 14272 14884 14278
rect 14752 14232 14832 14260
rect 14832 14214 14884 14220
rect 14844 12918 14872 14214
rect 15120 14074 15148 14282
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14916 13628 15292 13637
rect 14972 13626 14996 13628
rect 15052 13626 15076 13628
rect 15132 13626 15156 13628
rect 15212 13626 15236 13628
rect 14972 13574 14982 13626
rect 15226 13574 15236 13626
rect 14972 13572 14996 13574
rect 15052 13572 15076 13574
rect 15132 13572 15156 13574
rect 15212 13572 15236 13574
rect 14916 13563 15292 13572
rect 15396 13530 15424 14350
rect 15488 14278 15516 14470
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15396 12986 15424 13466
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14924 12776 14976 12782
rect 14752 12724 14924 12730
rect 14752 12718 14976 12724
rect 14752 12702 14964 12718
rect 14752 12306 14780 12702
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14752 11082 14780 12242
rect 14740 11076 14792 11082
rect 14740 11018 14792 11024
rect 14844 10674 14872 12582
rect 14916 12540 15292 12549
rect 14972 12538 14996 12540
rect 15052 12538 15076 12540
rect 15132 12538 15156 12540
rect 15212 12538 15236 12540
rect 14972 12486 14982 12538
rect 15226 12486 15236 12538
rect 14972 12484 14996 12486
rect 15052 12484 15076 12486
rect 15132 12484 15156 12486
rect 15212 12484 15236 12486
rect 14916 12475 15292 12484
rect 14916 11452 15292 11461
rect 14972 11450 14996 11452
rect 15052 11450 15076 11452
rect 15132 11450 15156 11452
rect 15212 11450 15236 11452
rect 14972 11398 14982 11450
rect 15226 11398 15236 11450
rect 14972 11396 14996 11398
rect 15052 11396 15076 11398
rect 15132 11396 15156 11398
rect 15212 11396 15236 11398
rect 14916 11387 15292 11396
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10742 15240 10950
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14476 10118 14596 10146
rect 13648 10084 13768 10112
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13544 10056 13596 10062
rect 13740 10044 13768 10084
rect 13820 10056 13872 10062
rect 13740 10016 13820 10044
rect 13544 9998 13596 10004
rect 14280 10056 14332 10062
rect 13820 9998 13872 10004
rect 14278 10024 14280 10033
rect 14332 10024 14334 10033
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13280 7970 13308 8842
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13372 8090 13400 8434
rect 13464 8294 13492 9454
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13280 7942 13400 7970
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13280 7546 13308 7822
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13372 6458 13400 7942
rect 13464 7342 13492 8230
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13556 6730 13584 9998
rect 13636 9988 13688 9994
rect 14278 9959 14334 9968
rect 13636 9930 13688 9936
rect 13648 8022 13676 9930
rect 14476 9602 14504 10118
rect 14660 10062 14688 10406
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14568 9722 14596 9998
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14372 9580 14424 9586
rect 14476 9574 14596 9602
rect 14372 9522 14424 9528
rect 14200 9178 14228 9522
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8634 13860 8774
rect 14384 8634 14412 9522
rect 14568 8838 14596 9574
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8634 14596 8774
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13648 7546 13676 7958
rect 13740 7546 13768 7958
rect 14384 7886 14412 8570
rect 14554 8528 14610 8537
rect 14554 8463 14556 8472
rect 14608 8463 14610 8472
rect 14556 8434 14608 8440
rect 14568 8362 14596 8434
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14188 7812 14240 7818
rect 14108 7772 14188 7800
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13740 6458 13768 7482
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13556 5642 13584 6190
rect 13740 5710 13768 6394
rect 14016 5710 14044 7346
rect 14108 7206 14136 7772
rect 14188 7754 14240 7760
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14568 7546 14596 7754
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14660 7002 14688 8026
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 11656 5468 12032 5477
rect 11712 5466 11736 5468
rect 11792 5466 11816 5468
rect 11872 5466 11896 5468
rect 11952 5466 11976 5468
rect 11712 5414 11722 5466
rect 11966 5414 11976 5466
rect 11712 5412 11736 5414
rect 11792 5412 11816 5414
rect 11872 5412 11896 5414
rect 11952 5412 11976 5414
rect 11656 5403 12032 5412
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4554 13032 4966
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11656 4380 12032 4389
rect 11712 4378 11736 4380
rect 11792 4378 11816 4380
rect 11872 4378 11896 4380
rect 11952 4378 11976 4380
rect 11712 4326 11722 4378
rect 11966 4326 11976 4378
rect 11712 4324 11736 4326
rect 11792 4324 11816 4326
rect 11872 4324 11896 4326
rect 11952 4324 11976 4326
rect 11656 4315 12032 4324
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 10916 3836 11292 3845
rect 10972 3834 10996 3836
rect 11052 3834 11076 3836
rect 11132 3834 11156 3836
rect 11212 3834 11236 3836
rect 10972 3782 10982 3834
rect 11226 3782 11236 3834
rect 10972 3780 10996 3782
rect 11052 3780 11076 3782
rect 11132 3780 11156 3782
rect 11212 3780 11236 3782
rect 10916 3771 11292 3780
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 11348 3466 11376 4014
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 11656 3292 12032 3301
rect 11712 3290 11736 3292
rect 11792 3290 11816 3292
rect 11872 3290 11896 3292
rect 11952 3290 11976 3292
rect 11712 3238 11722 3290
rect 11966 3238 11976 3290
rect 11712 3236 11736 3238
rect 11792 3236 11816 3238
rect 11872 3236 11896 3238
rect 11952 3236 11976 3238
rect 11656 3227 12032 3236
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 12084 3126 12112 3538
rect 12452 3534 12480 3878
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12268 3126 12296 3334
rect 13096 3126 13124 5102
rect 13188 4282 13216 5170
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13280 4214 13308 5238
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13648 4622 13676 5170
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13740 4146 13768 5646
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14108 5370 14136 5510
rect 14476 5370 14504 5510
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13832 4570 13860 4694
rect 14476 4622 14504 5306
rect 14660 4622 14688 6938
rect 14752 4826 14780 10542
rect 14844 10130 14872 10610
rect 14916 10364 15292 10373
rect 14972 10362 14996 10364
rect 15052 10362 15076 10364
rect 15132 10362 15156 10364
rect 15212 10362 15236 10364
rect 14972 10310 14982 10362
rect 15226 10310 15236 10362
rect 14972 10308 14996 10310
rect 15052 10308 15076 10310
rect 15132 10308 15156 10310
rect 15212 10308 15236 10310
rect 14916 10299 15292 10308
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14844 8974 14872 10066
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9722 15332 9930
rect 15292 9716 15344 9722
rect 15580 9674 15608 15506
rect 15656 15260 16032 15269
rect 15712 15258 15736 15260
rect 15792 15258 15816 15260
rect 15872 15258 15896 15260
rect 15952 15258 15976 15260
rect 15712 15206 15722 15258
rect 15966 15206 15976 15258
rect 15712 15204 15736 15206
rect 15792 15204 15816 15206
rect 15872 15204 15896 15206
rect 15952 15204 15976 15206
rect 15656 15195 16032 15204
rect 15750 14512 15806 14521
rect 15750 14447 15806 14456
rect 15764 14414 15792 14447
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15656 14172 16032 14181
rect 15712 14170 15736 14172
rect 15792 14170 15816 14172
rect 15872 14170 15896 14172
rect 15952 14170 15976 14172
rect 15712 14118 15722 14170
rect 15966 14118 15976 14170
rect 15712 14116 15736 14118
rect 15792 14116 15816 14118
rect 15872 14116 15896 14118
rect 15952 14116 15976 14118
rect 15656 14107 16032 14116
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15764 13530 15792 13874
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15856 13326 15884 13670
rect 16132 13410 16160 15642
rect 16224 13530 16252 21422
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16132 13382 16252 13410
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15656 13084 16032 13093
rect 15712 13082 15736 13084
rect 15792 13082 15816 13084
rect 15872 13082 15896 13084
rect 15952 13082 15976 13084
rect 15712 13030 15722 13082
rect 15966 13030 15976 13082
rect 15712 13028 15736 13030
rect 15792 13028 15816 13030
rect 15872 13028 15896 13030
rect 15952 13028 15976 13030
rect 15656 13019 16032 13028
rect 15656 11996 16032 12005
rect 15712 11994 15736 11996
rect 15792 11994 15816 11996
rect 15872 11994 15896 11996
rect 15952 11994 15976 11996
rect 15712 11942 15722 11994
rect 15966 11942 15976 11994
rect 15712 11940 15736 11942
rect 15792 11940 15816 11942
rect 15872 11940 15896 11942
rect 15952 11940 15976 11942
rect 15656 11931 16032 11940
rect 15656 10908 16032 10917
rect 15712 10906 15736 10908
rect 15792 10906 15816 10908
rect 15872 10906 15896 10908
rect 15952 10906 15976 10908
rect 15712 10854 15722 10906
rect 15966 10854 15976 10906
rect 15712 10852 15736 10854
rect 15792 10852 15816 10854
rect 15872 10852 15896 10854
rect 15952 10852 15976 10854
rect 15656 10843 16032 10852
rect 16224 10010 16252 13382
rect 16316 11286 16344 21490
rect 16408 18358 16436 25638
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16500 22982 16528 25298
rect 16684 23730 16712 25978
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 17236 23798 17264 25774
rect 17328 25158 17356 25978
rect 17420 25294 17448 26726
rect 17512 25906 17540 26794
rect 17604 26518 17632 26930
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17696 26450 17724 27406
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17696 26042 17724 26386
rect 17684 26036 17736 26042
rect 17684 25978 17736 25984
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17696 24993 17724 25842
rect 17880 25770 17908 26726
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17868 25764 17920 25770
rect 17868 25706 17920 25712
rect 17880 25430 17908 25706
rect 17972 25498 18000 26250
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 18064 26042 18092 26182
rect 18616 26042 18644 26930
rect 18052 26036 18104 26042
rect 18052 25978 18104 25984
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17868 25424 17920 25430
rect 17868 25366 17920 25372
rect 18064 25362 18092 25842
rect 18236 25764 18288 25770
rect 18236 25706 18288 25712
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 17682 24984 17738 24993
rect 18064 24954 18092 25298
rect 17682 24919 17738 24928
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 16948 23792 17000 23798
rect 16948 23734 17000 23740
rect 17224 23792 17276 23798
rect 17224 23734 17276 23740
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16684 23186 16712 23666
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16592 22545 16620 22918
rect 16684 22710 16712 23122
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16578 22536 16634 22545
rect 16578 22471 16634 22480
rect 16776 22030 16804 23462
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16960 21026 16988 23734
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17328 22642 17356 23258
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17316 22094 17368 22098
rect 17420 22094 17448 23054
rect 17972 22710 18000 23734
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17684 22568 17736 22574
rect 17684 22510 17736 22516
rect 17316 22092 17448 22094
rect 17368 22066 17448 22092
rect 17316 22034 17368 22040
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 16960 20998 17080 21026
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16500 19718 16528 20470
rect 16960 20398 16988 20878
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16960 19922 16988 20334
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16316 10810 16344 11018
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16316 10146 16344 10746
rect 16408 10266 16436 18158
rect 16500 17134 16528 19654
rect 16776 19446 16804 19790
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16868 18290 16896 18566
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17678 16804 18158
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17134 16804 17614
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16500 16794 16528 17070
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16500 15706 16528 16730
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16592 16017 16620 16594
rect 16684 16114 16712 16934
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16250 16804 16390
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16868 16114 16896 18226
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16578 16008 16634 16017
rect 16578 15943 16634 15952
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16868 15162 16896 15914
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16960 14414 16988 19314
rect 17052 18970 17080 20998
rect 17144 20942 17172 21898
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17052 18154 17080 18906
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 17052 16182 17080 16458
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17144 15978 17172 17206
rect 17236 16114 17264 17818
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17328 16250 17356 16390
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16500 14074 16528 14350
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16684 13326 16712 14350
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16500 12986 16528 13262
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16684 12434 16712 13262
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16776 12918 16804 13126
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16500 12406 16712 12434
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16316 10118 16436 10146
rect 16408 10062 16436 10118
rect 16132 9982 16252 10010
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16500 9994 16528 12406
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 9988 16540 9994
rect 15656 9820 16032 9829
rect 15712 9818 15736 9820
rect 15792 9818 15816 9820
rect 15872 9818 15896 9820
rect 15952 9818 15976 9820
rect 15712 9766 15722 9818
rect 15966 9766 15976 9818
rect 15712 9764 15736 9766
rect 15792 9764 15816 9766
rect 15872 9764 15896 9766
rect 15952 9764 15976 9766
rect 15656 9755 16032 9764
rect 15292 9658 15344 9664
rect 15396 9646 15608 9674
rect 14916 9276 15292 9285
rect 14972 9274 14996 9276
rect 15052 9274 15076 9276
rect 15132 9274 15156 9276
rect 15212 9274 15236 9276
rect 14972 9222 14982 9274
rect 15226 9222 15236 9274
rect 14972 9220 14996 9222
rect 15052 9220 15076 9222
rect 15132 9220 15156 9222
rect 15212 9220 15236 9222
rect 14916 9211 15292 9220
rect 15396 8974 15424 9646
rect 16132 9568 16160 9982
rect 16488 9930 16540 9936
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16224 9722 16252 9862
rect 16500 9738 16528 9930
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16316 9710 16528 9738
rect 16132 9540 16252 9568
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 14844 8566 14872 8910
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14916 8188 15292 8197
rect 14972 8186 14996 8188
rect 15052 8186 15076 8188
rect 15132 8186 15156 8188
rect 15212 8186 15236 8188
rect 14972 8134 14982 8186
rect 15226 8134 15236 8186
rect 14972 8132 14996 8134
rect 15052 8132 15076 8134
rect 15132 8132 15156 8134
rect 15212 8132 15236 8134
rect 14916 8123 15292 8132
rect 15396 7857 15424 8910
rect 15656 8732 16032 8741
rect 15712 8730 15736 8732
rect 15792 8730 15816 8732
rect 15872 8730 15896 8732
rect 15952 8730 15976 8732
rect 15712 8678 15722 8730
rect 15966 8678 15976 8730
rect 15712 8676 15736 8678
rect 15792 8676 15816 8678
rect 15872 8676 15896 8678
rect 15952 8676 15976 8678
rect 15656 8667 16032 8676
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 7886 15516 8230
rect 15476 7880 15528 7886
rect 15382 7848 15438 7857
rect 14832 7812 14884 7818
rect 15476 7822 15528 7828
rect 15382 7783 15438 7792
rect 14832 7754 14884 7760
rect 14844 7410 14872 7754
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14844 6798 14872 7346
rect 14916 7100 15292 7109
rect 14972 7098 14996 7100
rect 15052 7098 15076 7100
rect 15132 7098 15156 7100
rect 15212 7098 15236 7100
rect 14972 7046 14982 7098
rect 15226 7046 15236 7098
rect 14972 7044 14996 7046
rect 15052 7044 15076 7046
rect 15132 7044 15156 7046
rect 15212 7044 15236 7046
rect 14916 7035 15292 7044
rect 15396 7002 15424 7686
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15580 6798 15608 8298
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 8090 15700 8230
rect 15764 8090 15792 8434
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 15656 7644 16032 7653
rect 15712 7642 15736 7644
rect 15792 7642 15816 7644
rect 15872 7642 15896 7644
rect 15952 7642 15976 7644
rect 15712 7590 15722 7642
rect 15966 7590 15976 7642
rect 15712 7588 15736 7590
rect 15792 7588 15816 7590
rect 15872 7588 15896 7590
rect 15952 7588 15976 7590
rect 15656 7579 16032 7588
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 14844 5166 14872 6734
rect 15656 6556 16032 6565
rect 15712 6554 15736 6556
rect 15792 6554 15816 6556
rect 15872 6554 15896 6556
rect 15952 6554 15976 6556
rect 15712 6502 15722 6554
rect 15966 6502 15976 6554
rect 15712 6500 15736 6502
rect 15792 6500 15816 6502
rect 15872 6500 15896 6502
rect 15952 6500 15976 6502
rect 15656 6491 16032 6500
rect 14916 6012 15292 6021
rect 14972 6010 14996 6012
rect 15052 6010 15076 6012
rect 15132 6010 15156 6012
rect 15212 6010 15236 6012
rect 14972 5958 14982 6010
rect 15226 5958 15236 6010
rect 14972 5956 14996 5958
rect 15052 5956 15076 5958
rect 15132 5956 15156 5958
rect 15212 5956 15236 5958
rect 14916 5947 15292 5956
rect 15656 5468 16032 5477
rect 15712 5466 15736 5468
rect 15792 5466 15816 5468
rect 15872 5466 15896 5468
rect 15952 5466 15976 5468
rect 15712 5414 15722 5466
rect 15966 5414 15976 5466
rect 15712 5412 15736 5414
rect 15792 5412 15816 5414
rect 15872 5412 15896 5414
rect 15952 5412 15976 5414
rect 15656 5403 16032 5412
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14096 4616 14148 4622
rect 13832 4554 13952 4570
rect 14096 4558 14148 4564
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 13832 4548 13964 4554
rect 13832 4542 13912 4548
rect 13832 4282 13860 4542
rect 13912 4490 13964 4496
rect 14108 4282 14136 4558
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13280 3194 13308 3470
rect 13372 3194 13400 4082
rect 13740 3602 13768 4082
rect 14200 3738 14228 4082
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13740 3058 13768 3538
rect 14200 3194 14228 3674
rect 14476 3534 14504 4082
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 6916 2748 7292 2757
rect 6972 2746 6996 2748
rect 7052 2746 7076 2748
rect 7132 2746 7156 2748
rect 7212 2746 7236 2748
rect 6972 2694 6982 2746
rect 7226 2694 7236 2746
rect 6972 2692 6996 2694
rect 7052 2692 7076 2694
rect 7132 2692 7156 2694
rect 7212 2692 7236 2694
rect 6916 2683 7292 2692
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 8404 2582 8432 2994
rect 13740 2774 13768 2994
rect 14752 2854 14780 3538
rect 14844 3534 14872 5102
rect 14916 4924 15292 4933
rect 14972 4922 14996 4924
rect 15052 4922 15076 4924
rect 15132 4922 15156 4924
rect 15212 4922 15236 4924
rect 14972 4870 14982 4922
rect 15226 4870 15236 4922
rect 14972 4868 14996 4870
rect 15052 4868 15076 4870
rect 15132 4868 15156 4870
rect 15212 4868 15236 4870
rect 14916 4859 15292 4868
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14936 4078 14964 4626
rect 15656 4380 16032 4389
rect 15712 4378 15736 4380
rect 15792 4378 15816 4380
rect 15872 4378 15896 4380
rect 15952 4378 15976 4380
rect 15712 4326 15722 4378
rect 15966 4326 15976 4378
rect 15712 4324 15736 4326
rect 15792 4324 15816 4326
rect 15872 4324 15896 4326
rect 15952 4324 15976 4326
rect 15656 4315 16032 4324
rect 16132 4282 16160 7890
rect 16224 7750 16252 9540
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16224 5914 16252 6394
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16224 5778 16252 5850
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 16132 4026 16160 4218
rect 16316 4214 16344 9710
rect 16592 9602 16620 10202
rect 16684 10062 16712 11698
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16500 9574 16620 9602
rect 16408 8498 16436 9522
rect 16500 9110 16528 9574
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16500 8838 16528 9046
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16408 7954 16436 8434
rect 16592 7954 16620 8842
rect 16776 7970 16804 10746
rect 16868 9518 16896 13738
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16960 13326 16988 13670
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 17236 10554 17264 16050
rect 17420 16046 17448 22066
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 17604 20942 17632 21898
rect 17696 21894 17724 22510
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17880 21962 17908 22170
rect 18064 22094 18092 22986
rect 17972 22066 18092 22094
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17972 21690 18000 22066
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17604 19854 17632 20878
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17604 19718 17632 19790
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 18834 17632 19654
rect 17788 19378 17816 19790
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17512 18272 17540 18634
rect 17592 18284 17644 18290
rect 17512 18244 17592 18272
rect 17592 18226 17644 18232
rect 17604 18193 17632 18226
rect 17590 18184 17646 18193
rect 17590 18119 17646 18128
rect 17696 17882 17724 18634
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17512 17202 17540 17478
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17696 16658 17724 17070
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17604 14414 17632 16526
rect 17788 16289 17816 18090
rect 17880 18086 17908 20334
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17972 17678 18000 21626
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 18156 20398 18184 20810
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 19922 18184 20334
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17972 16674 18000 17614
rect 17880 16646 18000 16674
rect 17774 16280 17830 16289
rect 17774 16215 17830 16224
rect 17880 16130 17908 16646
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17972 16250 18000 16458
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17880 16102 18000 16130
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17880 15366 17908 15982
rect 17972 15366 18000 16102
rect 18064 15434 18092 19450
rect 18156 18834 18184 19858
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18156 18358 18184 18770
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18144 18148 18196 18154
rect 18144 18090 18196 18096
rect 18156 17116 18184 18090
rect 18248 17218 18276 25706
rect 18708 25294 18736 27270
rect 19444 27130 19472 27406
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19536 27062 19564 27406
rect 19656 27228 20032 27237
rect 19712 27226 19736 27228
rect 19792 27226 19816 27228
rect 19872 27226 19896 27228
rect 19952 27226 19976 27228
rect 19712 27174 19722 27226
rect 19966 27174 19976 27226
rect 19712 27172 19736 27174
rect 19792 27172 19816 27174
rect 19872 27172 19896 27174
rect 19952 27172 19976 27174
rect 19656 27163 20032 27172
rect 19524 27056 19576 27062
rect 19524 26998 19576 27004
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18800 26364 18828 26862
rect 20088 26790 20116 27406
rect 20352 27056 20404 27062
rect 20352 26998 20404 27004
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 18916 26684 19292 26693
rect 18972 26682 18996 26684
rect 19052 26682 19076 26684
rect 19132 26682 19156 26684
rect 19212 26682 19236 26684
rect 18972 26630 18982 26682
rect 19226 26630 19236 26682
rect 18972 26628 18996 26630
rect 19052 26628 19076 26630
rect 19132 26628 19156 26630
rect 19212 26628 19236 26630
rect 18916 26619 19292 26628
rect 18880 26376 18932 26382
rect 18800 26336 18880 26364
rect 18880 26318 18932 26324
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 18916 25596 19292 25605
rect 18972 25594 18996 25596
rect 19052 25594 19076 25596
rect 19132 25594 19156 25596
rect 19212 25594 19236 25596
rect 18972 25542 18982 25594
rect 19226 25542 19236 25594
rect 18972 25540 18996 25542
rect 19052 25540 19076 25542
rect 19132 25540 19156 25542
rect 19212 25540 19236 25542
rect 18916 25531 19292 25540
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 19352 24818 19380 25638
rect 19536 25498 19564 26250
rect 19656 26140 20032 26149
rect 19712 26138 19736 26140
rect 19792 26138 19816 26140
rect 19872 26138 19896 26140
rect 19952 26138 19976 26140
rect 19712 26086 19722 26138
rect 19966 26086 19976 26138
rect 19712 26084 19736 26086
rect 19792 26084 19816 26086
rect 19872 26084 19896 26086
rect 19952 26084 19976 26086
rect 19656 26075 20032 26084
rect 20088 26042 20116 26726
rect 20272 26314 20300 26726
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19656 25052 20032 25061
rect 19712 25050 19736 25052
rect 19792 25050 19816 25052
rect 19872 25050 19896 25052
rect 19952 25050 19976 25052
rect 19712 24998 19722 25050
rect 19966 24998 19976 25050
rect 19712 24996 19736 24998
rect 19792 24996 19816 24998
rect 19872 24996 19896 24998
rect 19952 24996 19976 24998
rect 19656 24987 20032 24996
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 18916 24508 19292 24517
rect 18972 24506 18996 24508
rect 19052 24506 19076 24508
rect 19132 24506 19156 24508
rect 19212 24506 19236 24508
rect 18972 24454 18982 24506
rect 19226 24454 19236 24506
rect 18972 24452 18996 24454
rect 19052 24452 19076 24454
rect 19132 24452 19156 24454
rect 19212 24452 19236 24454
rect 18916 24443 19292 24452
rect 19352 23882 19380 24754
rect 19536 24614 19564 24754
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19260 23854 19380 23882
rect 19260 23798 19288 23854
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 18340 23118 18368 23598
rect 18432 23526 18460 23666
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 18432 23186 18460 23462
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18340 21962 18368 23054
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18340 20942 18368 21898
rect 18432 21418 18460 22986
rect 18524 22030 18552 23462
rect 18916 23420 19292 23429
rect 18972 23418 18996 23420
rect 19052 23418 19076 23420
rect 19132 23418 19156 23420
rect 19212 23418 19236 23420
rect 18972 23366 18982 23418
rect 19226 23366 19236 23418
rect 18972 23364 18996 23366
rect 19052 23364 19076 23366
rect 19132 23364 19156 23366
rect 19212 23364 19236 23366
rect 18916 23355 19292 23364
rect 19444 23118 19472 23462
rect 19536 23254 19564 24550
rect 19904 24206 19932 24686
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 19656 23964 20032 23973
rect 19712 23962 19736 23964
rect 19792 23962 19816 23964
rect 19872 23962 19896 23964
rect 19952 23962 19976 23964
rect 19712 23910 19722 23962
rect 19966 23910 19976 23962
rect 19712 23908 19736 23910
rect 19792 23908 19816 23910
rect 19872 23908 19896 23910
rect 19952 23908 19976 23910
rect 19656 23899 20032 23908
rect 20088 23866 20116 24142
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 19524 23248 19576 23254
rect 19524 23190 19576 23196
rect 19432 23112 19484 23118
rect 19720 23100 19748 23734
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19812 23202 19840 23462
rect 19904 23322 19932 23666
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19984 23248 20036 23254
rect 19812 23174 19932 23202
rect 20036 23208 20116 23236
rect 19984 23190 20036 23196
rect 19904 23118 19932 23174
rect 19800 23112 19852 23118
rect 19432 23054 19484 23060
rect 19536 23072 19800 23100
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 18984 22710 19012 22986
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22710 19472 22918
rect 18972 22704 19024 22710
rect 18972 22646 19024 22652
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 18916 22332 19292 22341
rect 18972 22330 18996 22332
rect 19052 22330 19076 22332
rect 19132 22330 19156 22332
rect 19212 22330 19236 22332
rect 18972 22278 18982 22330
rect 19226 22278 19236 22330
rect 18972 22276 18996 22278
rect 19052 22276 19076 22278
rect 19132 22276 19156 22278
rect 19212 22276 19236 22278
rect 18916 22267 19292 22276
rect 19536 22234 19564 23072
rect 19892 23112 19944 23118
rect 19800 23054 19852 23060
rect 19890 23080 19892 23089
rect 19944 23080 19946 23089
rect 19890 23015 19946 23024
rect 19656 22876 20032 22885
rect 19712 22874 19736 22876
rect 19792 22874 19816 22876
rect 19872 22874 19896 22876
rect 19952 22874 19976 22876
rect 19712 22822 19722 22874
rect 19966 22822 19976 22874
rect 19712 22820 19736 22822
rect 19792 22820 19816 22822
rect 19872 22820 19896 22822
rect 19952 22820 19976 22822
rect 19656 22811 20032 22820
rect 20088 22710 20116 23208
rect 20180 22778 20208 24142
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20272 23662 20300 24006
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 20364 23066 20392 26998
rect 20548 26450 20576 27406
rect 21088 27328 21140 27334
rect 21088 27270 21140 27276
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 20548 25226 20576 26386
rect 20824 25226 20852 26930
rect 20916 26382 20944 27066
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20548 23186 20576 23666
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20272 23038 20392 23066
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 20076 22704 20128 22710
rect 19890 22672 19946 22681
rect 20076 22646 20128 22652
rect 19890 22607 19946 22616
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 19904 22137 19932 22607
rect 20088 22234 20116 22646
rect 20168 22636 20220 22642
rect 20272 22624 20300 23038
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20220 22596 20300 22624
rect 20168 22578 20220 22584
rect 20364 22522 20392 22918
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20180 22494 20392 22522
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19890 22128 19946 22137
rect 19248 22092 19300 22098
rect 19890 22063 19946 22072
rect 19248 22034 19300 22040
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18420 21412 18472 21418
rect 18420 21354 18472 21360
rect 18524 21078 18552 21966
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18512 21072 18564 21078
rect 18432 21020 18512 21026
rect 18432 21014 18564 21020
rect 18432 20998 18552 21014
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18340 20534 18368 20878
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18432 20398 18460 20998
rect 18616 20942 18644 21422
rect 18604 20936 18656 20942
rect 18524 20896 18604 20924
rect 18524 20466 18552 20896
rect 18604 20878 18656 20884
rect 18708 20806 18736 21966
rect 19260 21690 19288 22034
rect 19904 22030 19932 22063
rect 20088 22030 20116 22170
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 19524 21888 19576 21894
rect 19524 21830 19576 21836
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 18916 21244 19292 21253
rect 18972 21242 18996 21244
rect 19052 21242 19076 21244
rect 19132 21242 19156 21244
rect 19212 21242 19236 21244
rect 18972 21190 18982 21242
rect 19226 21190 19236 21242
rect 18972 21188 18996 21190
rect 19052 21188 19076 21190
rect 19132 21188 19156 21190
rect 19212 21188 19236 21190
rect 18916 21179 19292 21188
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18328 20392 18380 20398
rect 18326 20360 18328 20369
rect 18420 20392 18472 20398
rect 18380 20360 18382 20369
rect 18420 20334 18472 20340
rect 18326 20295 18382 20304
rect 18432 19786 18460 20334
rect 18524 19854 18552 20402
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18340 17626 18368 19722
rect 18432 19446 18460 19722
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 18432 18290 18460 19382
rect 18616 19378 18644 20538
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18616 18766 18644 19314
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18616 18222 18644 18702
rect 18708 18698 18736 20402
rect 18800 20262 18828 20810
rect 19340 20460 19392 20466
rect 19444 20448 19472 20946
rect 19536 20874 19564 21830
rect 19656 21788 20032 21797
rect 19712 21786 19736 21788
rect 19792 21786 19816 21788
rect 19872 21786 19896 21788
rect 19952 21786 19976 21788
rect 19712 21734 19722 21786
rect 19966 21734 19976 21786
rect 19712 21732 19736 21734
rect 19792 21732 19816 21734
rect 19872 21732 19896 21734
rect 19952 21732 19976 21734
rect 19656 21723 20032 21732
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19628 21146 19656 21626
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19628 20913 19656 21082
rect 19614 20904 19670 20913
rect 19524 20868 19576 20874
rect 19614 20839 19670 20848
rect 19524 20810 19576 20816
rect 19536 20534 19564 20810
rect 19656 20700 20032 20709
rect 19712 20698 19736 20700
rect 19792 20698 19816 20700
rect 19872 20698 19896 20700
rect 19952 20698 19976 20700
rect 19712 20646 19722 20698
rect 19966 20646 19976 20698
rect 19712 20644 19736 20646
rect 19792 20644 19816 20646
rect 19872 20644 19896 20646
rect 19952 20644 19976 20646
rect 19656 20635 20032 20644
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19392 20420 19472 20448
rect 19340 20402 19392 20408
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18340 17598 18552 17626
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18248 17190 18368 17218
rect 18156 17088 18276 17116
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 15910 18184 16390
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18052 15428 18104 15434
rect 18052 15370 18104 15376
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 18064 15178 18092 15370
rect 17696 15150 18092 15178
rect 17696 14890 17724 15150
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17328 10810 17356 13738
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17314 10704 17370 10713
rect 17314 10639 17316 10648
rect 17368 10639 17370 10648
rect 17316 10610 17368 10616
rect 17236 10526 17356 10554
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 16960 10062 16988 10406
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 9722 17080 9998
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16684 7942 16804 7970
rect 16500 7800 16528 7890
rect 16408 7772 16528 7800
rect 16580 7812 16632 7818
rect 16408 7274 16436 7772
rect 16580 7754 16632 7760
rect 16592 7698 16620 7754
rect 16500 7670 16620 7698
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16408 6254 16436 7210
rect 16500 7002 16528 7670
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16408 5370 16436 5510
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16408 4554 16436 5306
rect 16592 4622 16620 6666
rect 16684 5642 16712 7942
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16776 7546 16804 7822
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16868 5846 16896 9454
rect 17144 8090 17172 9522
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16868 5658 16896 5782
rect 17144 5778 17172 7482
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16776 5630 16896 5658
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16132 4010 16252 4026
rect 16132 4004 16264 4010
rect 16132 3998 16212 4004
rect 16212 3946 16264 3952
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 14916 3836 15292 3845
rect 14972 3834 14996 3836
rect 15052 3834 15076 3836
rect 15132 3834 15156 3836
rect 15212 3834 15236 3836
rect 14972 3782 14982 3834
rect 15226 3782 15236 3834
rect 14972 3780 14996 3782
rect 15052 3780 15076 3782
rect 15132 3780 15156 3782
rect 15212 3780 15236 3782
rect 14916 3771 15292 3780
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15396 3194 15424 3402
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15580 3058 15608 3878
rect 15656 3292 16032 3301
rect 15712 3290 15736 3292
rect 15792 3290 15816 3292
rect 15872 3290 15896 3292
rect 15952 3290 15976 3292
rect 15712 3238 15722 3290
rect 15966 3238 15976 3290
rect 15712 3236 15736 3238
rect 15792 3236 15816 3238
rect 15872 3236 15896 3238
rect 15952 3236 15976 3238
rect 15656 3227 16032 3236
rect 16132 3058 16160 3878
rect 16224 3398 16252 3946
rect 16408 3738 16436 4082
rect 16684 4078 16712 5578
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16776 3738 16804 5630
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16868 5234 16896 5510
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17236 4826 17264 10406
rect 17328 9674 17356 10526
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 10266 17448 10406
rect 17498 10296 17554 10305
rect 17408 10260 17460 10266
rect 17498 10231 17500 10240
rect 17408 10202 17460 10208
rect 17552 10231 17554 10240
rect 17500 10202 17552 10208
rect 17604 10112 17632 14350
rect 17696 10674 17724 14826
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17696 10130 17724 10610
rect 17512 10084 17632 10112
rect 17684 10124 17736 10130
rect 17408 10056 17460 10062
rect 17512 10044 17540 10084
rect 17684 10066 17736 10072
rect 17460 10016 17540 10044
rect 17590 10024 17646 10033
rect 17408 9998 17460 10004
rect 17590 9959 17646 9968
rect 17328 9646 17540 9674
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17420 9178 17448 9522
rect 17512 9382 17540 9646
rect 17604 9586 17632 9959
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17328 7342 17356 8910
rect 17420 8634 17448 9114
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17328 5234 17356 7278
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17328 4282 17356 4558
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17420 4146 17448 4490
rect 17512 4146 17540 9318
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17604 7546 17632 8026
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17788 7342 17816 11154
rect 17880 10266 17908 15030
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18064 13326 18092 13942
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 12986 18092 13262
rect 18156 13258 18184 15846
rect 18248 15473 18276 17088
rect 18234 15464 18290 15473
rect 18234 15399 18290 15408
rect 18248 13394 18276 15399
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17880 8634 17908 9522
rect 17972 8922 18000 12650
rect 18064 9586 18092 12718
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 9178 18092 9318
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17972 8894 18092 8922
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17972 7154 18000 8774
rect 17788 7126 18000 7154
rect 17788 6390 17816 7126
rect 18064 6882 18092 8894
rect 17972 6854 18092 6882
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 4282 17908 4422
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 17880 4146 17908 4218
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17420 3738 17448 4082
rect 17972 3942 18000 6854
rect 18050 6760 18106 6769
rect 18050 6695 18106 6704
rect 18064 5710 18092 6695
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18156 4282 18184 13194
rect 18248 12782 18276 13330
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18248 9654 18276 10950
rect 18340 10146 18368 17190
rect 18432 16794 18460 17478
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18524 16538 18552 17598
rect 18616 17105 18644 17682
rect 18602 17096 18658 17105
rect 18602 17031 18658 17040
rect 18432 16510 18552 16538
rect 18432 16454 18460 16510
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 16250 18552 16390
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18432 15162 18460 15982
rect 18524 15502 18552 16186
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18616 15094 18644 17031
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18708 14550 18736 16594
rect 18800 16590 18828 20198
rect 18916 20156 19292 20165
rect 18972 20154 18996 20156
rect 19052 20154 19076 20156
rect 19132 20154 19156 20156
rect 19212 20154 19236 20156
rect 18972 20102 18982 20154
rect 19226 20102 19236 20154
rect 18972 20100 18996 20102
rect 19052 20100 19076 20102
rect 19132 20100 19156 20102
rect 19212 20100 19236 20102
rect 18916 20091 19292 20100
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18984 19378 19012 19858
rect 19536 19854 19564 20198
rect 19628 19922 19656 20470
rect 19892 20460 19944 20466
rect 20088 20448 20116 21966
rect 20180 21350 20208 22494
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20364 21554 20392 22374
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20180 20466 20208 21286
rect 20272 20942 20300 21354
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 19944 20420 20116 20448
rect 20168 20460 20220 20466
rect 19892 20402 19944 20408
rect 20168 20402 20220 20408
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19720 19922 19748 20334
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19812 19854 19840 20334
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19800 19848 19852 19854
rect 19904 19836 19932 20402
rect 20076 19848 20128 19854
rect 19904 19808 20076 19836
rect 19800 19790 19852 19796
rect 20076 19790 20128 19796
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18916 19068 19292 19077
rect 18972 19066 18996 19068
rect 19052 19066 19076 19068
rect 19132 19066 19156 19068
rect 19212 19066 19236 19068
rect 18972 19014 18982 19066
rect 19226 19014 19236 19066
rect 18972 19012 18996 19014
rect 19052 19012 19076 19014
rect 19132 19012 19156 19014
rect 19212 19012 19236 19014
rect 18916 19003 19292 19012
rect 19352 18834 19380 19722
rect 19812 19700 19840 19790
rect 19536 19672 19840 19700
rect 19536 19378 19564 19672
rect 19656 19612 20032 19621
rect 19712 19610 19736 19612
rect 19792 19610 19816 19612
rect 19872 19610 19896 19612
rect 19952 19610 19976 19612
rect 19712 19558 19722 19610
rect 19966 19558 19976 19610
rect 19712 19556 19736 19558
rect 19792 19556 19816 19558
rect 19872 19556 19896 19558
rect 19952 19556 19976 19558
rect 19656 19547 20032 19556
rect 20088 19378 20116 19790
rect 20180 19514 20208 20402
rect 20272 20058 20300 20538
rect 20364 20398 20392 21490
rect 20456 21468 20484 22578
rect 20548 22506 20576 23122
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 20534 21992 20590 22001
rect 20534 21927 20590 21936
rect 20548 21622 20576 21927
rect 20536 21616 20588 21622
rect 20536 21558 20588 21564
rect 20536 21480 20588 21486
rect 20456 21440 20536 21468
rect 20536 21422 20588 21428
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20456 20534 20484 20742
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20272 19718 20300 19994
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19536 19174 19564 19314
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18892 18358 18920 18634
rect 19720 18630 19748 19314
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19656 18524 20032 18533
rect 19712 18522 19736 18524
rect 19792 18522 19816 18524
rect 19872 18522 19896 18524
rect 19952 18522 19976 18524
rect 19712 18470 19722 18522
rect 19966 18470 19976 18522
rect 19712 18468 19736 18470
rect 19792 18468 19816 18470
rect 19872 18468 19896 18470
rect 19952 18468 19976 18470
rect 19656 18459 20032 18468
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18916 17980 19292 17989
rect 18972 17978 18996 17980
rect 19052 17978 19076 17980
rect 19132 17978 19156 17980
rect 19212 17978 19236 17980
rect 18972 17926 18982 17978
rect 19226 17926 19236 17978
rect 18972 17924 18996 17926
rect 19052 17924 19076 17926
rect 19132 17924 19156 17926
rect 19212 17924 19236 17926
rect 18916 17915 19292 17924
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 16980 19288 17614
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19352 17338 19380 17546
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19352 17082 19380 17274
rect 19444 17270 19472 17478
rect 19656 17436 20032 17445
rect 19712 17434 19736 17436
rect 19792 17434 19816 17436
rect 19872 17434 19896 17436
rect 19952 17434 19976 17436
rect 19712 17382 19722 17434
rect 19966 17382 19976 17434
rect 19712 17380 19736 17382
rect 19792 17380 19816 17382
rect 19872 17380 19896 17382
rect 19952 17380 19976 17382
rect 19656 17371 20032 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19352 17054 19564 17082
rect 19432 16992 19484 16998
rect 19260 16952 19380 16980
rect 18916 16892 19292 16901
rect 18972 16890 18996 16892
rect 19052 16890 19076 16892
rect 19132 16890 19156 16892
rect 19212 16890 19236 16892
rect 18972 16838 18982 16890
rect 19226 16838 19236 16890
rect 18972 16836 18996 16838
rect 19052 16836 19076 16838
rect 19132 16836 19156 16838
rect 19212 16836 19236 16838
rect 18916 16827 19292 16836
rect 19248 16788 19300 16794
rect 19352 16776 19380 16952
rect 19432 16934 19484 16940
rect 19300 16748 19380 16776
rect 19248 16730 19300 16736
rect 19444 16590 19472 16934
rect 18788 16584 18840 16590
rect 19248 16584 19300 16590
rect 18788 16526 18840 16532
rect 18970 16552 19026 16561
rect 19248 16526 19300 16532
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 18970 16487 19026 16496
rect 18786 16280 18842 16289
rect 18984 16250 19012 16487
rect 18786 16215 18842 16224
rect 18972 16244 19024 16250
rect 18800 16182 18828 16215
rect 18972 16186 19024 16192
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 19260 16114 19288 16526
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19338 16280 19394 16289
rect 19338 16215 19340 16224
rect 19392 16215 19394 16224
rect 19340 16186 19392 16192
rect 19352 16114 19380 16186
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18800 14618 18828 15982
rect 18916 15804 19292 15813
rect 18972 15802 18996 15804
rect 19052 15802 19076 15804
rect 19132 15802 19156 15804
rect 19212 15802 19236 15804
rect 18972 15750 18982 15802
rect 19226 15750 19236 15802
rect 18972 15748 18996 15750
rect 19052 15748 19076 15750
rect 19132 15748 19156 15750
rect 19212 15748 19236 15750
rect 18916 15739 19292 15748
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19352 15162 19380 15574
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 18916 14716 19292 14725
rect 18972 14714 18996 14716
rect 19052 14714 19076 14716
rect 19132 14714 19156 14716
rect 19212 14714 19236 14716
rect 18972 14662 18982 14714
rect 19226 14662 19236 14714
rect 18972 14660 18996 14662
rect 19052 14660 19076 14662
rect 19132 14660 19156 14662
rect 19212 14660 19236 14662
rect 18916 14651 19292 14660
rect 19352 14618 19380 14962
rect 19444 14618 19472 16390
rect 19536 16114 19564 17054
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19616 16720 19668 16726
rect 19616 16662 19668 16668
rect 19628 16454 19656 16662
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19656 16348 20032 16357
rect 19712 16346 19736 16348
rect 19792 16346 19816 16348
rect 19872 16346 19896 16348
rect 19952 16346 19976 16348
rect 19712 16294 19722 16346
rect 19966 16294 19976 16346
rect 19712 16292 19736 16294
rect 19792 16292 19816 16294
rect 19872 16292 19896 16294
rect 19952 16292 19976 16294
rect 19656 16283 20032 16292
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 20088 15706 20116 16730
rect 20180 16114 20208 19246
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 19656 15260 20032 15269
rect 19712 15258 19736 15260
rect 19792 15258 19816 15260
rect 19872 15258 19896 15260
rect 19952 15258 19976 15260
rect 19712 15206 19722 15258
rect 19966 15206 19976 15258
rect 19712 15204 19736 15206
rect 19792 15204 19816 15206
rect 19872 15204 19896 15206
rect 19952 15204 19976 15206
rect 19656 15195 20032 15204
rect 20088 15162 20116 15370
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18696 14408 18748 14414
rect 18694 14376 18696 14385
rect 18880 14408 18932 14414
rect 18748 14376 18750 14385
rect 18604 14340 18656 14346
rect 18880 14350 18932 14356
rect 18694 14311 18750 14320
rect 18604 14282 18656 14288
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18432 13530 18460 13738
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18432 13433 18460 13466
rect 18616 13462 18644 14282
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18604 13456 18656 13462
rect 18418 13424 18474 13433
rect 18604 13398 18656 13404
rect 18418 13359 18474 13368
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12986 18552 13126
rect 18708 12986 18736 13942
rect 18800 13530 18828 14214
rect 18892 14074 18920 14350
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 19352 13870 19380 14554
rect 19444 13938 19472 14554
rect 19656 14172 20032 14181
rect 19712 14170 19736 14172
rect 19792 14170 19816 14172
rect 19872 14170 19896 14172
rect 19952 14170 19976 14172
rect 19712 14118 19722 14170
rect 19966 14118 19976 14170
rect 19712 14116 19736 14118
rect 19792 14116 19816 14118
rect 19872 14116 19896 14118
rect 19952 14116 19976 14118
rect 19656 14107 20032 14116
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19340 13864 19392 13870
rect 19392 13812 19472 13818
rect 19340 13806 19472 13812
rect 19352 13790 19472 13806
rect 18916 13628 19292 13637
rect 18972 13626 18996 13628
rect 19052 13626 19076 13628
rect 19132 13626 19156 13628
rect 19212 13626 19236 13628
rect 18972 13574 18982 13626
rect 19226 13574 19236 13626
rect 18972 13572 18996 13574
rect 19052 13572 19076 13574
rect 19132 13572 19156 13574
rect 19212 13572 19236 13574
rect 18916 13563 19292 13572
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19260 12986 19288 13398
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18800 12238 18828 12582
rect 18916 12540 19292 12549
rect 18972 12538 18996 12540
rect 19052 12538 19076 12540
rect 19132 12538 19156 12540
rect 19212 12538 19236 12540
rect 18972 12486 18982 12538
rect 19226 12486 19236 12538
rect 18972 12484 18996 12486
rect 19052 12484 19076 12486
rect 19132 12484 19156 12486
rect 19212 12484 19236 12486
rect 18916 12475 19292 12484
rect 19352 12442 19380 13194
rect 19444 12986 19472 13790
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19536 12918 19564 13670
rect 19656 13084 20032 13093
rect 19712 13082 19736 13084
rect 19792 13082 19816 13084
rect 19872 13082 19896 13084
rect 19952 13082 19976 13084
rect 19712 13030 19722 13082
rect 19966 13030 19976 13082
rect 19712 13028 19736 13030
rect 19792 13028 19816 13030
rect 19872 13028 19896 13030
rect 19952 13028 19976 13030
rect 19656 13019 20032 13028
rect 20088 12986 20116 13874
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18916 11452 19292 11461
rect 18972 11450 18996 11452
rect 19052 11450 19076 11452
rect 19132 11450 19156 11452
rect 19212 11450 19236 11452
rect 18972 11398 18982 11450
rect 19226 11398 19236 11450
rect 18972 11396 18996 11398
rect 19052 11396 19076 11398
rect 19132 11396 19156 11398
rect 19212 11396 19236 11398
rect 18916 11387 19292 11396
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10810 18460 10950
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18602 10296 18658 10305
rect 18602 10231 18658 10240
rect 18340 10118 18552 10146
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18248 8090 18276 9590
rect 18340 9042 18368 9998
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9722 18460 9862
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18432 7562 18460 9522
rect 18340 7534 18460 7562
rect 18340 4690 18368 7534
rect 18524 7478 18552 10118
rect 18616 8294 18644 10231
rect 18708 9450 18736 11086
rect 18880 11008 18932 11014
rect 18800 10968 18880 10996
rect 18800 9994 18828 10968
rect 18880 10950 18932 10956
rect 18916 10364 19292 10373
rect 18972 10362 18996 10364
rect 19052 10362 19076 10364
rect 19132 10362 19156 10364
rect 19212 10362 19236 10364
rect 18972 10310 18982 10362
rect 19226 10310 19236 10362
rect 18972 10308 18996 10310
rect 19052 10308 19076 10310
rect 19132 10308 19156 10310
rect 19212 10308 19236 10310
rect 18916 10299 19292 10308
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18892 9364 18920 10202
rect 19444 9674 19472 12718
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 19656 11996 20032 12005
rect 19712 11994 19736 11996
rect 19792 11994 19816 11996
rect 19872 11994 19896 11996
rect 19952 11994 19976 11996
rect 19712 11942 19722 11994
rect 19966 11942 19976 11994
rect 19712 11940 19736 11942
rect 19792 11940 19816 11942
rect 19872 11940 19896 11942
rect 19952 11940 19976 11942
rect 19656 11931 20032 11940
rect 20180 11830 20208 12038
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19536 10674 19564 11222
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 19656 10908 20032 10917
rect 19712 10906 19736 10908
rect 19792 10906 19816 10908
rect 19872 10906 19896 10908
rect 19952 10906 19976 10908
rect 19712 10854 19722 10906
rect 19966 10854 19976 10906
rect 19712 10852 19736 10854
rect 19792 10852 19816 10854
rect 19872 10852 19896 10854
rect 19952 10852 19976 10854
rect 19656 10843 20032 10852
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 20180 10554 20208 11018
rect 20272 10742 20300 19654
rect 20364 19378 20392 19858
rect 20456 19786 20484 20470
rect 20548 20262 20576 21422
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20640 16810 20668 25094
rect 20824 23118 20852 25162
rect 20916 23594 20944 26318
rect 20904 23588 20956 23594
rect 20904 23530 20956 23536
rect 20916 23236 20944 23530
rect 20916 23208 21036 23236
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20720 22568 20772 22574
rect 20824 22556 20852 23054
rect 20772 22528 20852 22556
rect 20720 22510 20772 22516
rect 20916 22166 20944 23054
rect 21008 22982 21036 23208
rect 21100 23050 21128 27270
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 21088 23044 21140 23050
rect 21088 22986 21140 22992
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 21100 22642 21128 22986
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21192 22506 21220 25298
rect 21180 22500 21232 22506
rect 21180 22442 21232 22448
rect 20904 22160 20956 22166
rect 20718 22128 20774 22137
rect 20904 22102 20956 22108
rect 20718 22063 20774 22072
rect 20732 20466 20760 22063
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20824 21350 20852 21830
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20916 20398 20944 22102
rect 21284 21690 21312 26318
rect 21640 26240 21692 26246
rect 21640 26182 21692 26188
rect 21364 25832 21416 25838
rect 21364 25774 21416 25780
rect 21376 24750 21404 25774
rect 21652 25362 21680 26182
rect 22112 25974 22140 26318
rect 22100 25968 22152 25974
rect 22100 25910 22152 25916
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 21192 19514 21220 21490
rect 21376 21418 21404 24006
rect 22112 23798 22140 25774
rect 22480 25430 22508 25774
rect 22468 25424 22520 25430
rect 22468 25366 22520 25372
rect 22572 25294 22600 29315
rect 22916 27772 23292 27781
rect 22972 27770 22996 27772
rect 23052 27770 23076 27772
rect 23132 27770 23156 27772
rect 23212 27770 23236 27772
rect 22972 27718 22982 27770
rect 23226 27718 23236 27770
rect 22972 27716 22996 27718
rect 23052 27716 23076 27718
rect 23132 27716 23156 27718
rect 23212 27716 23236 27718
rect 22916 27707 23292 27716
rect 23656 27228 24032 27237
rect 23712 27226 23736 27228
rect 23792 27226 23816 27228
rect 23872 27226 23896 27228
rect 23952 27226 23976 27228
rect 23712 27174 23722 27226
rect 23966 27174 23976 27226
rect 23712 27172 23736 27174
rect 23792 27172 23816 27174
rect 23872 27172 23896 27174
rect 23952 27172 23976 27174
rect 23656 27163 24032 27172
rect 22916 26684 23292 26693
rect 22972 26682 22996 26684
rect 23052 26682 23076 26684
rect 23132 26682 23156 26684
rect 23212 26682 23236 26684
rect 22972 26630 22982 26682
rect 23226 26630 23236 26682
rect 22972 26628 22996 26630
rect 23052 26628 23076 26630
rect 23132 26628 23156 26630
rect 23212 26628 23236 26630
rect 22916 26619 23292 26628
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22664 25158 22692 25978
rect 23492 25974 23520 26250
rect 23656 26140 24032 26149
rect 23712 26138 23736 26140
rect 23792 26138 23816 26140
rect 23872 26138 23896 26140
rect 23952 26138 23976 26140
rect 23712 26086 23722 26138
rect 23966 26086 23976 26138
rect 23712 26084 23736 26086
rect 23792 26084 23816 26086
rect 23872 26084 23896 26086
rect 23952 26084 23976 26086
rect 23656 26075 24032 26084
rect 23480 25968 23532 25974
rect 23480 25910 23532 25916
rect 23572 25764 23624 25770
rect 23572 25706 23624 25712
rect 22916 25596 23292 25605
rect 22972 25594 22996 25596
rect 23052 25594 23076 25596
rect 23132 25594 23156 25596
rect 23212 25594 23236 25596
rect 22972 25542 22982 25594
rect 23226 25542 23236 25594
rect 22972 25540 22996 25542
rect 23052 25540 23076 25542
rect 23132 25540 23156 25542
rect 23212 25540 23236 25542
rect 22916 25531 23292 25540
rect 23584 25362 23612 25706
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22664 24206 22692 25094
rect 22916 24508 23292 24517
rect 22972 24506 22996 24508
rect 23052 24506 23076 24508
rect 23132 24506 23156 24508
rect 23212 24506 23236 24508
rect 22972 24454 22982 24506
rect 23226 24454 23236 24506
rect 22972 24452 22996 24454
rect 23052 24452 23076 24454
rect 23132 24452 23156 24454
rect 23212 24452 23236 24454
rect 22916 24443 23292 24452
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22100 23792 22152 23798
rect 22100 23734 22152 23740
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21744 22642 21772 23258
rect 22112 23186 22140 23734
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22388 23254 22416 23598
rect 22376 23248 22428 23254
rect 22376 23190 22428 23196
rect 22664 23202 22692 24142
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22848 23662 22876 24074
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23216 23730 23244 24006
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 23388 23656 23440 23662
rect 23388 23598 23440 23604
rect 22916 23420 23292 23429
rect 22972 23418 22996 23420
rect 23052 23418 23076 23420
rect 23132 23418 23156 23420
rect 23212 23418 23236 23420
rect 22972 23366 22982 23418
rect 23226 23366 23236 23418
rect 22972 23364 22996 23366
rect 23052 23364 23076 23366
rect 23132 23364 23156 23366
rect 23212 23364 23236 23366
rect 22916 23355 23292 23364
rect 22664 23186 22784 23202
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 22664 23180 22796 23186
rect 22664 23174 22744 23180
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21560 22030 21588 22510
rect 21744 22030 21772 22578
rect 21916 22500 21968 22506
rect 21916 22442 21968 22448
rect 21928 22166 21956 22442
rect 21916 22160 21968 22166
rect 21916 22102 21968 22108
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21744 21690 21772 21966
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21364 21412 21416 21418
rect 21364 21354 21416 21360
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21928 19786 21956 21286
rect 22112 21078 22140 23122
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 22204 22778 22232 23054
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22296 22234 22324 22510
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22204 21622 22232 21966
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22664 21554 22692 23174
rect 22744 23122 22796 23128
rect 23400 22642 23428 23598
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23492 22506 23520 24210
rect 23584 23526 23612 25298
rect 23656 25052 24032 25061
rect 23712 25050 23736 25052
rect 23792 25050 23816 25052
rect 23872 25050 23896 25052
rect 23952 25050 23976 25052
rect 23712 24998 23722 25050
rect 23966 24998 23976 25050
rect 23712 24996 23736 24998
rect 23792 24996 23816 24998
rect 23872 24996 23896 24998
rect 23952 24996 23976 24998
rect 23656 24987 24032 24996
rect 24504 24993 24532 29315
rect 24490 24984 24546 24993
rect 24490 24919 24546 24928
rect 25136 24132 25188 24138
rect 25136 24074 25188 24080
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 23656 23964 24032 23973
rect 23712 23962 23736 23964
rect 23792 23962 23816 23964
rect 23872 23962 23896 23964
rect 23952 23962 23976 23964
rect 23712 23910 23722 23962
rect 23966 23910 23976 23962
rect 23712 23908 23736 23910
rect 23792 23908 23816 23910
rect 23872 23908 23896 23910
rect 23952 23908 23976 23910
rect 23656 23899 24032 23908
rect 24504 23798 24532 24006
rect 24492 23792 24544 23798
rect 24492 23734 24544 23740
rect 25148 23526 25176 24074
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 23584 22658 23612 23462
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 23656 22876 24032 22885
rect 23712 22874 23736 22876
rect 23792 22874 23816 22876
rect 23872 22874 23896 22876
rect 23952 22874 23976 22876
rect 23712 22822 23722 22874
rect 23966 22822 23976 22874
rect 23712 22820 23736 22822
rect 23792 22820 23816 22822
rect 23872 22820 23896 22822
rect 23952 22820 23976 22822
rect 23656 22811 24032 22820
rect 24228 22710 24256 22918
rect 24504 22710 24532 22918
rect 24216 22704 24268 22710
rect 23584 22630 23704 22658
rect 24216 22646 24268 22652
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 23480 22500 23532 22506
rect 23480 22442 23532 22448
rect 22916 22332 23292 22341
rect 22972 22330 22996 22332
rect 23052 22330 23076 22332
rect 23132 22330 23156 22332
rect 23212 22330 23236 22332
rect 22972 22278 22982 22330
rect 23226 22278 23236 22330
rect 22972 22276 22996 22278
rect 23052 22276 23076 22278
rect 23132 22276 23156 22278
rect 23212 22276 23236 22278
rect 22916 22267 23292 22276
rect 23492 22166 23520 22442
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23676 22094 23704 22630
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 23952 22234 23980 22510
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23584 22066 23704 22094
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22100 21072 22152 21078
rect 22100 21014 22152 21020
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 22020 19922 22048 20198
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22112 19786 22140 21014
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 20398 22232 20742
rect 22664 20466 22692 21490
rect 23492 21486 23520 21830
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 22916 21244 23292 21253
rect 22972 21242 22996 21244
rect 23052 21242 23076 21244
rect 23132 21242 23156 21244
rect 23212 21242 23236 21244
rect 22972 21190 22982 21242
rect 23226 21190 23236 21242
rect 22972 21188 22996 21190
rect 23052 21188 23076 21190
rect 23132 21188 23156 21190
rect 23212 21188 23236 21190
rect 22916 21179 23292 21188
rect 23584 21162 23612 22066
rect 24124 21956 24176 21962
rect 24124 21898 24176 21904
rect 23656 21788 24032 21797
rect 23712 21786 23736 21788
rect 23792 21786 23816 21788
rect 23872 21786 23896 21788
rect 23952 21786 23976 21788
rect 23712 21734 23722 21786
rect 23966 21734 23976 21786
rect 23712 21732 23736 21734
rect 23792 21732 23816 21734
rect 23872 21732 23896 21734
rect 23952 21732 23976 21734
rect 23656 21723 24032 21732
rect 24136 21486 24164 21898
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24228 21350 24256 22646
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24412 21690 24440 21966
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 23492 21134 23612 21162
rect 23492 20942 23520 21134
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22192 20392 22244 20398
rect 22192 20334 22244 20340
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 21916 19780 21968 19786
rect 21916 19722 21968 19728
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 22112 19174 22140 19722
rect 22480 19514 22508 19858
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22112 18290 22140 19110
rect 22204 18970 22232 19314
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22572 18766 22600 20334
rect 23492 20262 23520 20878
rect 24228 20874 24256 21286
rect 24216 20868 24268 20874
rect 24216 20810 24268 20816
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 22916 20156 23292 20165
rect 22972 20154 22996 20156
rect 23052 20154 23076 20156
rect 23132 20154 23156 20156
rect 23212 20154 23236 20156
rect 22972 20102 22982 20154
rect 23226 20102 23236 20154
rect 22972 20100 22996 20102
rect 23052 20100 23076 20102
rect 23132 20100 23156 20102
rect 23212 20100 23236 20102
rect 22916 20091 23292 20100
rect 23584 20058 23612 20742
rect 23656 20700 24032 20709
rect 23712 20698 23736 20700
rect 23792 20698 23816 20700
rect 23872 20698 23896 20700
rect 23952 20698 23976 20700
rect 23712 20646 23722 20698
rect 23966 20646 23976 20698
rect 23712 20644 23736 20646
rect 23792 20644 23816 20646
rect 23872 20644 23896 20646
rect 23952 20644 23976 20646
rect 23656 20635 24032 20644
rect 24136 20534 24164 20742
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23676 19768 23704 20198
rect 24136 19854 24164 20334
rect 24124 19848 24176 19854
rect 24124 19790 24176 19796
rect 23584 19740 23704 19768
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22112 17882 22140 18226
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 20456 16782 20668 16810
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20364 16250 20392 16526
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20456 15978 20484 16782
rect 20628 16720 20680 16726
rect 20628 16662 20680 16668
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20548 16182 20576 16390
rect 20536 16176 20588 16182
rect 20536 16118 20588 16124
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20444 14884 20496 14890
rect 20444 14826 20496 14832
rect 20456 11082 20484 14826
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20180 10526 20300 10554
rect 19656 9820 20032 9829
rect 19712 9818 19736 9820
rect 19792 9818 19816 9820
rect 19872 9818 19896 9820
rect 19952 9818 19976 9820
rect 19712 9766 19722 9818
rect 19966 9766 19976 9818
rect 19712 9764 19736 9766
rect 19792 9764 19816 9766
rect 19872 9764 19896 9766
rect 19952 9764 19976 9766
rect 19656 9755 20032 9764
rect 19352 9646 19472 9674
rect 19352 9518 19380 9646
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 18800 9336 18920 9364
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18432 5370 18460 7414
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 10916 2748 11292 2757
rect 10972 2746 10996 2748
rect 11052 2746 11076 2748
rect 11132 2746 11156 2748
rect 11212 2746 11236 2748
rect 10972 2694 10982 2746
rect 11226 2694 11236 2746
rect 10972 2692 10996 2694
rect 11052 2692 11076 2694
rect 11132 2692 11156 2694
rect 11212 2692 11236 2694
rect 10916 2683 11292 2692
rect 13648 2746 13768 2774
rect 14916 2748 15292 2757
rect 14972 2746 14996 2748
rect 15052 2746 15076 2748
rect 15132 2746 15156 2748
rect 15212 2746 15236 2748
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 13648 2514 13676 2746
rect 14972 2694 14982 2746
rect 15226 2694 15236 2746
rect 14972 2692 14996 2694
rect 15052 2692 15076 2694
rect 15132 2692 15156 2694
rect 15212 2692 15236 2694
rect 14916 2683 15292 2692
rect 16224 2582 16252 3334
rect 16316 3194 16344 3402
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 17972 3126 18000 3878
rect 18340 3398 18368 4014
rect 18432 3602 18460 5306
rect 18524 4758 18552 6734
rect 18616 6322 18644 7346
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18708 6304 18736 7278
rect 18800 7206 18828 9336
rect 18916 9276 19292 9285
rect 18972 9274 18996 9276
rect 19052 9274 19076 9276
rect 19132 9274 19156 9276
rect 19212 9274 19236 9276
rect 18972 9222 18982 9274
rect 19226 9222 19236 9274
rect 18972 9220 18996 9222
rect 19052 9220 19076 9222
rect 19132 9220 19156 9222
rect 19212 9220 19236 9222
rect 18916 9211 19292 9220
rect 18916 8188 19292 8197
rect 18972 8186 18996 8188
rect 19052 8186 19076 8188
rect 19132 8186 19156 8188
rect 19212 8186 19236 8188
rect 18972 8134 18982 8186
rect 19226 8134 19236 8186
rect 18972 8132 18996 8134
rect 19052 8132 19076 8134
rect 19132 8132 19156 8134
rect 19212 8132 19236 8134
rect 18916 8123 19292 8132
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18916 7100 19292 7109
rect 18972 7098 18996 7100
rect 19052 7098 19076 7100
rect 19132 7098 19156 7100
rect 19212 7098 19236 7100
rect 18972 7046 18982 7098
rect 19226 7046 19236 7098
rect 18972 7044 18996 7046
rect 19052 7044 19076 7046
rect 19132 7044 19156 7046
rect 19212 7044 19236 7046
rect 18916 7035 19292 7044
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18800 6458 18828 6938
rect 19352 6882 19380 9454
rect 19656 8732 20032 8741
rect 19712 8730 19736 8732
rect 19792 8730 19816 8732
rect 19872 8730 19896 8732
rect 19952 8730 19976 8732
rect 19712 8678 19722 8730
rect 19966 8678 19976 8730
rect 19712 8676 19736 8678
rect 19792 8676 19816 8678
rect 19872 8676 19896 8678
rect 19952 8676 19976 8678
rect 19656 8667 20032 8676
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 19444 7886 19472 8366
rect 19708 8016 19760 8022
rect 19706 7984 19708 7993
rect 19760 7984 19762 7993
rect 19706 7919 19762 7928
rect 19812 7886 19840 8366
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19800 7880 19852 7886
rect 19996 7868 20024 8366
rect 20180 8022 20208 8366
rect 20168 8016 20220 8022
rect 20168 7958 20220 7964
rect 20076 7880 20128 7886
rect 19996 7840 20076 7868
rect 19800 7822 19852 7828
rect 20076 7822 20128 7828
rect 19444 7546 19472 7822
rect 19524 7812 19576 7818
rect 19524 7754 19576 7760
rect 19432 7540 19484 7546
rect 19536 7528 19564 7754
rect 19656 7644 20032 7653
rect 19712 7642 19736 7644
rect 19792 7642 19816 7644
rect 19872 7642 19896 7644
rect 19952 7642 19976 7644
rect 19712 7590 19722 7642
rect 19966 7590 19976 7642
rect 19712 7588 19736 7590
rect 19792 7588 19816 7590
rect 19872 7588 19896 7590
rect 19952 7588 19976 7590
rect 19656 7579 20032 7588
rect 19536 7500 19840 7528
rect 19432 7482 19484 7488
rect 19168 6854 19380 6882
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18788 6316 18840 6322
rect 18708 6276 18788 6304
rect 18616 5642 18644 6258
rect 18708 5846 18736 6276
rect 18788 6258 18840 6264
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5636 18656 5642
rect 18604 5578 18656 5584
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18524 4010 18552 4694
rect 18616 4146 18644 5578
rect 18708 5234 18736 5782
rect 18800 5710 18828 6122
rect 19168 6118 19196 6854
rect 19444 6730 19472 7482
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19536 7002 19564 7346
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19260 6186 19288 6666
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 18916 6012 19292 6021
rect 18972 6010 18996 6012
rect 19052 6010 19076 6012
rect 19132 6010 19156 6012
rect 19212 6010 19236 6012
rect 18972 5958 18982 6010
rect 19226 5958 19236 6010
rect 18972 5956 18996 5958
rect 19052 5956 19076 5958
rect 19132 5956 19156 5958
rect 19212 5956 19236 5958
rect 18916 5947 19292 5956
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18708 4214 18736 5170
rect 18800 5098 18828 5646
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 18984 5234 19012 5578
rect 19352 5386 19380 6598
rect 19444 6322 19472 6666
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19444 5914 19472 6054
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19536 5778 19564 6938
rect 19720 6798 19748 7278
rect 19812 6798 19840 7500
rect 20088 7410 20116 7822
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19656 6556 20032 6565
rect 19712 6554 19736 6556
rect 19792 6554 19816 6556
rect 19872 6554 19896 6556
rect 19952 6554 19976 6556
rect 19712 6502 19722 6554
rect 19966 6502 19976 6554
rect 19712 6500 19736 6502
rect 19792 6500 19816 6502
rect 19872 6500 19896 6502
rect 19952 6500 19976 6502
rect 19656 6491 20032 6500
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19352 5358 19472 5386
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18800 4554 18828 5034
rect 18916 4924 19292 4933
rect 18972 4922 18996 4924
rect 19052 4922 19076 4924
rect 19132 4922 19156 4924
rect 19212 4922 19236 4924
rect 18972 4870 18982 4922
rect 19226 4870 19236 4922
rect 18972 4868 18996 4870
rect 19052 4868 19076 4870
rect 19132 4868 19156 4870
rect 19212 4868 19236 4870
rect 18916 4859 19292 4868
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18916 3836 19292 3845
rect 18972 3834 18996 3836
rect 19052 3834 19076 3836
rect 19132 3834 19156 3836
rect 19212 3834 19236 3836
rect 18972 3782 18982 3834
rect 19226 3782 19236 3834
rect 18972 3780 18996 3782
rect 19052 3780 19076 3782
rect 19132 3780 19156 3782
rect 19212 3780 19236 3782
rect 18916 3771 19292 3780
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18340 3194 18368 3334
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18800 3126 18828 3334
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18916 2748 19292 2757
rect 18972 2746 18996 2748
rect 19052 2746 19076 2748
rect 19132 2746 19156 2748
rect 19212 2746 19236 2748
rect 18972 2694 18982 2746
rect 19226 2694 19236 2746
rect 18972 2692 18996 2694
rect 19052 2692 19076 2694
rect 19132 2692 19156 2694
rect 19212 2692 19236 2694
rect 18916 2683 19292 2692
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 3656 2204 4032 2213
rect 3712 2202 3736 2204
rect 3792 2202 3816 2204
rect 3872 2202 3896 2204
rect 3952 2202 3976 2204
rect 3712 2150 3722 2202
rect 3966 2150 3976 2202
rect 3712 2148 3736 2150
rect 3792 2148 3816 2150
rect 3872 2148 3896 2150
rect 3952 2148 3976 2150
rect 3656 2139 4032 2148
rect 5828 800 5856 2382
rect 7656 2204 8032 2213
rect 7712 2202 7736 2204
rect 7792 2202 7816 2204
rect 7872 2202 7896 2204
rect 7952 2202 7976 2204
rect 7712 2150 7722 2202
rect 7966 2150 7976 2202
rect 7712 2148 7736 2150
rect 7792 2148 7816 2150
rect 7872 2148 7896 2150
rect 7952 2148 7976 2150
rect 7656 2139 8032 2148
rect 8404 800 8432 2382
rect 11656 2204 12032 2213
rect 11712 2202 11736 2204
rect 11792 2202 11816 2204
rect 11872 2202 11896 2204
rect 11952 2202 11976 2204
rect 11712 2150 11722 2202
rect 11966 2150 11976 2202
rect 11712 2148 11736 2150
rect 11792 2148 11816 2150
rect 11872 2148 11896 2150
rect 11952 2148 11976 2150
rect 11656 2139 12032 2148
rect 12820 1306 12848 2382
rect 15656 2204 16032 2213
rect 15712 2202 15736 2204
rect 15792 2202 15816 2204
rect 15872 2202 15896 2204
rect 15952 2202 15976 2204
rect 15712 2150 15722 2202
rect 15966 2150 15976 2202
rect 15712 2148 15736 2150
rect 15792 2148 15816 2150
rect 15872 2148 15896 2150
rect 15952 2148 15976 2150
rect 15656 2139 16032 2148
rect 12820 1278 12940 1306
rect 12912 800 12940 1278
rect 16132 800 16160 2382
rect 19352 800 19380 5238
rect 19444 4622 19472 5358
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19536 4146 19564 5714
rect 19628 5710 19656 6054
rect 20088 5710 20116 7346
rect 20180 7342 20208 7958
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20272 6780 20300 10526
rect 20640 8650 20668 16662
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20732 13326 20760 13806
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 12306 20760 13262
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20824 11354 20852 12174
rect 21008 11898 21036 16594
rect 21468 16522 21496 16934
rect 21560 16658 21588 17070
rect 22112 16998 22140 17818
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22296 17626 22324 17682
rect 22204 17598 22324 17626
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22112 16794 22140 16934
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21560 16114 21588 16594
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21836 16182 21864 16390
rect 21824 16176 21876 16182
rect 21822 16144 21824 16153
rect 21876 16144 21878 16153
rect 21548 16108 21600 16114
rect 21822 16079 21878 16088
rect 21548 16050 21600 16056
rect 21560 15638 21588 16050
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21192 14482 21220 15574
rect 21836 15502 21864 15914
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 14958 21864 15438
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21836 13870 21864 14894
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22020 13394 22048 13806
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21192 12306 21220 12582
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 22020 11898 22048 12786
rect 22204 12442 22232 17598
rect 22480 17338 22508 18158
rect 22572 17746 22600 18702
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22572 17134 22600 17682
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22572 16182 22600 17070
rect 22664 16454 22692 19246
rect 22916 19068 23292 19077
rect 22972 19066 22996 19068
rect 23052 19066 23076 19068
rect 23132 19066 23156 19068
rect 23212 19066 23236 19068
rect 22972 19014 22982 19066
rect 23226 19014 23236 19066
rect 22972 19012 22996 19014
rect 23052 19012 23076 19014
rect 23132 19012 23156 19014
rect 23212 19012 23236 19014
rect 22916 19003 23292 19012
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23400 18426 23428 18702
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 22916 17980 23292 17989
rect 22972 17978 22996 17980
rect 23052 17978 23076 17980
rect 23132 17978 23156 17980
rect 23212 17978 23236 17980
rect 22972 17926 22982 17978
rect 23226 17926 23236 17978
rect 22972 17924 22996 17926
rect 23052 17924 23076 17926
rect 23132 17924 23156 17926
rect 23212 17924 23236 17926
rect 22916 17915 23292 17924
rect 23400 17746 23428 18362
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23492 17882 23520 18158
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 22836 17264 22888 17270
rect 22836 17206 22888 17212
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22848 16250 22876 17206
rect 22916 16892 23292 16901
rect 22972 16890 22996 16892
rect 23052 16890 23076 16892
rect 23132 16890 23156 16892
rect 23212 16890 23236 16892
rect 22972 16838 22982 16890
rect 23226 16838 23236 16890
rect 22972 16836 22996 16838
rect 23052 16836 23076 16838
rect 23132 16836 23156 16838
rect 23212 16836 23236 16838
rect 22916 16827 23292 16836
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22916 15804 23292 15813
rect 22972 15802 22996 15804
rect 23052 15802 23076 15804
rect 23132 15802 23156 15804
rect 23212 15802 23236 15804
rect 22972 15750 22982 15802
rect 23226 15750 23236 15802
rect 22972 15748 22996 15750
rect 23052 15748 23076 15750
rect 23132 15748 23156 15750
rect 23212 15748 23236 15750
rect 22916 15739 23292 15748
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22848 15094 22876 15302
rect 22836 15088 22888 15094
rect 22836 15030 22888 15036
rect 22916 14716 23292 14725
rect 22972 14714 22996 14716
rect 23052 14714 23076 14716
rect 23132 14714 23156 14716
rect 23212 14714 23236 14716
rect 22972 14662 22982 14714
rect 23226 14662 23236 14714
rect 22972 14660 22996 14662
rect 23052 14660 23076 14662
rect 23132 14660 23156 14662
rect 23212 14660 23236 14662
rect 22916 14651 23292 14660
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 14006 22324 14214
rect 22284 14000 22336 14006
rect 22284 13942 22336 13948
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22848 13530 22876 13942
rect 22916 13628 23292 13637
rect 22972 13626 22996 13628
rect 23052 13626 23076 13628
rect 23132 13626 23156 13628
rect 23212 13626 23236 13628
rect 22972 13574 22982 13626
rect 23226 13574 23236 13626
rect 22972 13572 22996 13574
rect 23052 13572 23076 13574
rect 23132 13572 23156 13574
rect 23212 13572 23236 13574
rect 22916 13563 23292 13572
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 22916 12540 23292 12549
rect 22972 12538 22996 12540
rect 23052 12538 23076 12540
rect 23132 12538 23156 12540
rect 23212 12538 23236 12540
rect 22972 12486 22982 12538
rect 23226 12486 23236 12538
rect 22972 12484 22996 12486
rect 23052 12484 23076 12486
rect 23132 12484 23156 12486
rect 23212 12484 23236 12486
rect 22916 12475 23292 12484
rect 22192 12436 22244 12442
rect 23400 12434 23428 17206
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23492 14414 23520 15438
rect 23584 14482 23612 19740
rect 23656 19612 24032 19621
rect 23712 19610 23736 19612
rect 23792 19610 23816 19612
rect 23872 19610 23896 19612
rect 23952 19610 23976 19612
rect 23712 19558 23722 19610
rect 23966 19558 23976 19610
rect 23712 19556 23736 19558
rect 23792 19556 23816 19558
rect 23872 19556 23896 19558
rect 23952 19556 23976 19558
rect 23656 19547 24032 19556
rect 23656 18524 24032 18533
rect 23712 18522 23736 18524
rect 23792 18522 23816 18524
rect 23872 18522 23896 18524
rect 23952 18522 23976 18524
rect 23712 18470 23722 18522
rect 23966 18470 23976 18522
rect 23712 18468 23736 18470
rect 23792 18468 23816 18470
rect 23872 18468 23896 18470
rect 23952 18468 23976 18470
rect 23656 18459 24032 18468
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23860 17882 23888 18294
rect 24136 18086 24164 19790
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23656 17436 24032 17445
rect 23712 17434 23736 17436
rect 23792 17434 23816 17436
rect 23872 17434 23896 17436
rect 23952 17434 23976 17436
rect 23712 17382 23722 17434
rect 23966 17382 23976 17434
rect 23712 17380 23736 17382
rect 23792 17380 23816 17382
rect 23872 17380 23896 17382
rect 23952 17380 23976 17382
rect 23656 17371 24032 17380
rect 23656 16348 24032 16357
rect 23712 16346 23736 16348
rect 23792 16346 23816 16348
rect 23872 16346 23896 16348
rect 23952 16346 23976 16348
rect 23712 16294 23722 16346
rect 23966 16294 23976 16346
rect 23712 16292 23736 16294
rect 23792 16292 23816 16294
rect 23872 16292 23896 16294
rect 23952 16292 23976 16294
rect 23656 16283 24032 16292
rect 23656 15260 24032 15269
rect 23712 15258 23736 15260
rect 23792 15258 23816 15260
rect 23872 15258 23896 15260
rect 23952 15258 23976 15260
rect 23712 15206 23722 15258
rect 23966 15206 23976 15258
rect 23712 15204 23736 15206
rect 23792 15204 23816 15206
rect 23872 15204 23896 15206
rect 23952 15204 23976 15206
rect 23656 15195 24032 15204
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 24136 14414 24164 14962
rect 24228 14958 24256 20810
rect 24412 20602 24440 21626
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24584 21480 24636 21486
rect 24584 21422 24636 21428
rect 24400 20596 24452 20602
rect 24400 20538 24452 20544
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24412 19990 24440 20198
rect 24400 19984 24452 19990
rect 24400 19926 24452 19932
rect 24400 16516 24452 16522
rect 24400 16458 24452 16464
rect 24412 15502 24440 16458
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24412 14414 24440 15438
rect 24596 15434 24624 21422
rect 24780 21146 24808 21490
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24780 20942 24808 21082
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24964 20602 24992 21286
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 24688 20058 24716 20334
rect 25148 20244 25176 23462
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25240 22098 25268 22578
rect 26514 22536 26570 22545
rect 26514 22471 26516 22480
rect 26568 22471 26570 22480
rect 26516 22442 26568 22448
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25424 21554 25452 22374
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25516 20466 25544 21286
rect 25700 20874 25728 21286
rect 25688 20868 25740 20874
rect 25688 20810 25740 20816
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25228 20256 25280 20262
rect 25148 20216 25228 20244
rect 25228 20198 25280 20204
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 25240 19854 25268 20198
rect 25516 19990 25544 20402
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 25792 19854 25820 20402
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25044 18692 25096 18698
rect 25044 18634 25096 18640
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24872 17882 24900 18294
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 24688 15026 24716 15506
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24688 14482 24716 14758
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 23656 14172 24032 14181
rect 23712 14170 23736 14172
rect 23792 14170 23816 14172
rect 23872 14170 23896 14172
rect 23952 14170 23976 14172
rect 23712 14118 23722 14170
rect 23966 14118 23976 14170
rect 23712 14116 23736 14118
rect 23792 14116 23816 14118
rect 23872 14116 23896 14118
rect 23952 14116 23976 14118
rect 23656 14107 24032 14116
rect 24136 13938 24164 14350
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 22192 12378 22244 12384
rect 22848 12406 23428 12434
rect 22204 11898 22232 12378
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11898 22784 12174
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 21008 11150 21036 11834
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21376 11218 21404 11562
rect 21468 11218 21496 11630
rect 21744 11354 21772 11766
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 21468 10606 21496 11154
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21468 10130 21496 10542
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21468 9042 21496 10066
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 20548 8634 20668 8650
rect 20536 8628 20668 8634
rect 20588 8622 20668 8628
rect 20536 8570 20588 8576
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20548 7886 20576 8298
rect 20640 8242 20668 8622
rect 20732 8537 20760 8842
rect 20718 8528 20774 8537
rect 20718 8463 20774 8472
rect 20732 8362 20760 8463
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20640 8214 20760 8242
rect 20732 8090 20760 8214
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20456 7410 20484 7754
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20456 7206 20484 7346
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20180 6752 20300 6780
rect 20180 6458 20208 6752
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20272 5710 20300 6394
rect 20364 5930 20392 7142
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20456 6254 20484 6938
rect 20548 6798 20576 7822
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20732 6866 20760 7278
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20548 6390 20576 6734
rect 20640 6390 20668 6734
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20548 6202 20576 6326
rect 20732 6322 20760 6802
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20548 6174 20760 6202
rect 20364 5902 20668 5930
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 19656 5468 20032 5477
rect 19712 5466 19736 5468
rect 19792 5466 19816 5468
rect 19872 5466 19896 5468
rect 19952 5466 19976 5468
rect 19712 5414 19722 5466
rect 19966 5414 19976 5466
rect 19712 5412 19736 5414
rect 19792 5412 19816 5414
rect 19872 5412 19896 5414
rect 19952 5412 19976 5414
rect 19656 5403 20032 5412
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19812 4622 19840 4762
rect 19996 4622 20024 5102
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19656 4380 20032 4389
rect 19712 4378 19736 4380
rect 19792 4378 19816 4380
rect 19872 4378 19896 4380
rect 19952 4378 19976 4380
rect 19712 4326 19722 4378
rect 19966 4326 19976 4378
rect 19712 4324 19736 4326
rect 19792 4324 19816 4326
rect 19872 4324 19896 4326
rect 19952 4324 19976 4326
rect 19656 4315 20032 4324
rect 20088 4282 20116 5646
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 20180 4162 20208 5034
rect 20272 4622 20300 5646
rect 20364 5234 20392 5782
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20456 5234 20484 5578
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20364 4826 20392 5170
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20548 4554 20576 4762
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 19996 4146 20208 4162
rect 20548 4146 20576 4490
rect 20640 4486 20668 5902
rect 20732 5234 20760 6174
rect 20824 6118 20852 7754
rect 21100 7342 21128 8366
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6934 20944 7142
rect 20904 6928 20956 6934
rect 20904 6870 20956 6876
rect 20916 6361 20944 6870
rect 20994 6760 21050 6769
rect 20994 6695 21050 6704
rect 21008 6662 21036 6695
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 20902 6352 20958 6361
rect 20902 6287 20958 6296
rect 20916 6186 20944 6287
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20824 5778 20852 6054
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20824 5234 20852 5714
rect 21100 5710 21128 7278
rect 21192 5846 21220 7822
rect 21284 7478 21312 8842
rect 21468 8498 21496 8978
rect 21560 8634 21588 11018
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21744 10130 21772 10406
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21928 9654 21956 10678
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21652 8498 21680 8910
rect 21928 8566 21956 9590
rect 22112 9382 22140 11086
rect 22480 9518 22508 11630
rect 22756 11150 22784 11834
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22848 9586 22876 12406
rect 23388 11688 23440 11694
rect 23388 11630 23440 11636
rect 22916 11452 23292 11461
rect 22972 11450 22996 11452
rect 23052 11450 23076 11452
rect 23132 11450 23156 11452
rect 23212 11450 23236 11452
rect 22972 11398 22982 11450
rect 23226 11398 23236 11450
rect 22972 11396 22996 11398
rect 23052 11396 23076 11398
rect 23132 11396 23156 11398
rect 23212 11396 23236 11398
rect 22916 11387 23292 11396
rect 23400 11218 23428 11630
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 22916 10364 23292 10373
rect 22972 10362 22996 10364
rect 23052 10362 23076 10364
rect 23132 10362 23156 10364
rect 23212 10362 23236 10364
rect 22972 10310 22982 10362
rect 23226 10310 23236 10362
rect 22972 10308 22996 10310
rect 23052 10308 23076 10310
rect 23132 10308 23156 10310
rect 23212 10308 23236 10310
rect 22916 10299 23292 10308
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21284 6934 21312 7414
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 21284 6798 21312 6870
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21376 6118 21404 8230
rect 21836 7954 21864 8366
rect 21928 7954 21956 8502
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21640 7880 21692 7886
rect 21692 7840 21772 7868
rect 21640 7822 21692 7828
rect 21744 7342 21772 7840
rect 21732 7336 21784 7342
rect 21638 7304 21694 7313
rect 21732 7278 21784 7284
rect 21638 7239 21640 7248
rect 21692 7239 21694 7248
rect 21640 7210 21692 7216
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21560 6390 21588 6666
rect 21652 6458 21680 6734
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21192 5710 21220 5782
rect 21744 5778 21772 6394
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21836 5710 21864 7890
rect 21928 7002 21956 7890
rect 22204 7886 22232 8230
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22480 7410 22508 7754
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22388 7274 22416 7346
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 21916 6996 21968 7002
rect 21916 6938 21968 6944
rect 21928 6322 21956 6938
rect 22112 6798 22140 7142
rect 22100 6792 22152 6798
rect 22152 6740 22324 6746
rect 22100 6734 22324 6740
rect 22112 6718 22324 6734
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22098 6352 22154 6361
rect 21916 6316 21968 6322
rect 22204 6322 22232 6598
rect 22296 6322 22324 6718
rect 22098 6287 22100 6296
rect 21916 6258 21968 6264
rect 22152 6287 22154 6296
rect 22192 6316 22244 6322
rect 22100 6258 22152 6264
rect 22192 6258 22244 6264
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22112 6202 22140 6258
rect 22112 6174 22232 6202
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20824 5098 20852 5170
rect 21008 5166 21036 5646
rect 21100 5302 21128 5646
rect 21088 5296 21140 5302
rect 21088 5238 21140 5244
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20812 5092 20864 5098
rect 20812 5034 20864 5040
rect 20824 4622 20852 5034
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20628 4480 20680 4486
rect 21008 4468 21036 5102
rect 21928 4622 21956 6054
rect 22112 4826 22140 6054
rect 22204 5710 22232 6174
rect 22296 5778 22324 6258
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22204 4622 22232 5510
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21088 4480 21140 4486
rect 21008 4440 21088 4468
rect 20628 4422 20680 4428
rect 21088 4422 21140 4428
rect 21100 4214 21128 4422
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19984 4140 20208 4146
rect 20036 4134 20208 4140
rect 20536 4140 20588 4146
rect 19984 4082 20036 4088
rect 20536 4082 20588 4088
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21468 3534 21496 3878
rect 21928 3738 21956 4558
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22112 4214 22140 4422
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22480 3942 22508 7346
rect 22572 6798 22600 8910
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22572 5710 22600 6598
rect 22664 6254 22692 9318
rect 22848 8498 22876 9522
rect 23308 9466 23336 9862
rect 23308 9438 23428 9466
rect 22916 9276 23292 9285
rect 22972 9274 22996 9276
rect 23052 9274 23076 9276
rect 23132 9274 23156 9276
rect 23212 9274 23236 9276
rect 22972 9222 22982 9274
rect 23226 9222 23236 9274
rect 22972 9220 22996 9222
rect 23052 9220 23076 9222
rect 23132 9220 23156 9222
rect 23212 9220 23236 9222
rect 22916 9211 23292 9220
rect 23400 9042 23428 9438
rect 23492 9330 23520 13806
rect 24136 13326 24164 13874
rect 24412 13870 24440 14350
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 23656 13084 24032 13093
rect 23712 13082 23736 13084
rect 23792 13082 23816 13084
rect 23872 13082 23896 13084
rect 23952 13082 23976 13084
rect 23712 13030 23722 13082
rect 23966 13030 23976 13082
rect 23712 13028 23736 13030
rect 23792 13028 23816 13030
rect 23872 13028 23896 13030
rect 23952 13028 23976 13030
rect 23656 13019 24032 13028
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23584 11830 23612 12038
rect 23656 11996 24032 12005
rect 23712 11994 23736 11996
rect 23792 11994 23816 11996
rect 23872 11994 23896 11996
rect 23952 11994 23976 11996
rect 23712 11942 23722 11994
rect 23966 11942 23976 11994
rect 23712 11940 23736 11942
rect 23792 11940 23816 11942
rect 23872 11940 23896 11942
rect 23952 11940 23976 11942
rect 23656 11931 24032 11940
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 24136 11082 24164 13262
rect 24412 12986 24440 13806
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 23656 10908 24032 10917
rect 23712 10906 23736 10908
rect 23792 10906 23816 10908
rect 23872 10906 23896 10908
rect 23952 10906 23976 10908
rect 23712 10854 23722 10906
rect 23966 10854 23976 10906
rect 23712 10852 23736 10854
rect 23792 10852 23816 10854
rect 23872 10852 23896 10854
rect 23952 10852 23976 10854
rect 23656 10843 24032 10852
rect 24136 10062 24164 11018
rect 24504 10810 24532 12038
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 23656 9820 24032 9829
rect 23712 9818 23736 9820
rect 23792 9818 23816 9820
rect 23872 9818 23896 9820
rect 23952 9818 23976 9820
rect 23712 9766 23722 9818
rect 23966 9766 23976 9818
rect 23712 9764 23736 9766
rect 23792 9764 23816 9766
rect 23872 9764 23896 9766
rect 23952 9764 23976 9766
rect 23656 9755 24032 9764
rect 24596 9586 24624 12582
rect 24780 12238 24808 17546
rect 25056 17338 25084 18634
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 11626 24808 12174
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24688 10810 24716 11018
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24872 10062 24900 14214
rect 24952 14000 25004 14006
rect 24952 13942 25004 13948
rect 24964 12850 24992 13942
rect 25056 13394 25084 15302
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 25148 14346 25176 14758
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25240 13734 25268 19790
rect 25792 18426 25820 19790
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 26068 18290 26096 21490
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 25964 18080 26016 18086
rect 25964 18022 26016 18028
rect 25976 17270 26004 18022
rect 26068 17678 26096 18226
rect 26160 17882 26188 20810
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26436 19718 26464 20334
rect 26424 19712 26476 19718
rect 26424 19654 26476 19660
rect 26436 18970 26464 19654
rect 26424 18964 26476 18970
rect 26424 18906 26476 18912
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 26252 18426 26280 18634
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 26068 17542 26096 17614
rect 26056 17536 26108 17542
rect 26056 17478 26108 17484
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25976 15434 26004 15846
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25228 13728 25280 13734
rect 25976 13705 26004 14894
rect 25228 13670 25280 13676
rect 25962 13696 26018 13705
rect 25962 13631 26018 13640
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 24952 12844 25004 12850
rect 24952 12786 25004 12792
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24964 11694 24992 12242
rect 25792 12238 25820 13126
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24964 10674 24992 11630
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25700 11082 25728 11494
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 25056 10062 25084 10678
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25148 10266 25176 10542
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 23940 9376 23992 9382
rect 23492 9302 23704 9330
rect 23940 9318 23992 9324
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23584 9058 23612 9114
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23492 9030 23612 9058
rect 23492 8906 23520 9030
rect 23676 8974 23704 9302
rect 23952 8974 23980 9318
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 23480 8900 23532 8906
rect 23480 8842 23532 8848
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22756 7410 22784 8230
rect 22848 7886 22876 8434
rect 22916 8188 23292 8197
rect 22972 8186 22996 8188
rect 23052 8186 23076 8188
rect 23132 8186 23156 8188
rect 23212 8186 23236 8188
rect 22972 8134 22982 8186
rect 23226 8134 23236 8186
rect 22972 8132 22996 8134
rect 23052 8132 23076 8134
rect 23132 8132 23156 8134
rect 23212 8132 23236 8134
rect 22916 8123 23292 8132
rect 23296 7948 23348 7954
rect 23348 7908 23428 7936
rect 23296 7890 23348 7896
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22756 7274 22784 7346
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22848 6882 22876 7822
rect 22916 7100 23292 7109
rect 22972 7098 22996 7100
rect 23052 7098 23076 7100
rect 23132 7098 23156 7100
rect 23212 7098 23236 7100
rect 22972 7046 22982 7098
rect 23226 7046 23236 7098
rect 22972 7044 22996 7046
rect 23052 7044 23076 7046
rect 23132 7044 23156 7046
rect 23212 7044 23236 7046
rect 22916 7035 23292 7044
rect 22756 6854 22876 6882
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22664 4622 22692 6190
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22572 4214 22600 4422
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 19656 3292 20032 3301
rect 19712 3290 19736 3292
rect 19792 3290 19816 3292
rect 19872 3290 19896 3292
rect 19952 3290 19976 3292
rect 19712 3238 19722 3290
rect 19966 3238 19976 3290
rect 19712 3236 19736 3238
rect 19792 3236 19816 3238
rect 19872 3236 19896 3238
rect 19952 3236 19976 3238
rect 19656 3227 20032 3236
rect 21468 2990 21496 3470
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22480 3194 22508 3402
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22664 3058 22692 4558
rect 22756 3602 22784 6854
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 22836 6724 22888 6730
rect 22836 6666 22888 6672
rect 22848 6322 22876 6666
rect 23124 6322 23152 6734
rect 23400 6458 23428 7908
rect 23492 7426 23520 8842
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23584 8090 23612 8774
rect 23656 8732 24032 8741
rect 23712 8730 23736 8732
rect 23792 8730 23816 8732
rect 23872 8730 23896 8732
rect 23952 8730 23976 8732
rect 23712 8678 23722 8730
rect 23966 8678 23976 8730
rect 23712 8676 23736 8678
rect 23792 8676 23816 8678
rect 23872 8676 23896 8678
rect 23952 8676 23976 8678
rect 23656 8667 24032 8676
rect 24136 8634 24164 8910
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24124 8424 24176 8430
rect 24228 8412 24256 9454
rect 24780 8974 24808 9998
rect 24872 9042 24900 9998
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9178 24992 9862
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24952 8900 25004 8906
rect 25056 8888 25084 9998
rect 25240 9586 25268 9998
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25136 9104 25188 9110
rect 25136 9046 25188 9052
rect 25004 8860 25084 8888
rect 24952 8842 25004 8848
rect 24176 8384 24256 8412
rect 24124 8366 24176 8372
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23656 7644 24032 7653
rect 23712 7642 23736 7644
rect 23792 7642 23816 7644
rect 23872 7642 23896 7644
rect 23952 7642 23976 7644
rect 23712 7590 23722 7642
rect 23966 7590 23976 7642
rect 23712 7588 23736 7590
rect 23792 7588 23816 7590
rect 23872 7588 23896 7590
rect 23952 7588 23976 7590
rect 23656 7579 24032 7588
rect 23492 7410 23612 7426
rect 23492 7404 23624 7410
rect 23492 7398 23572 7404
rect 23572 7346 23624 7352
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23584 6458 23612 6734
rect 23656 6556 24032 6565
rect 23712 6554 23736 6556
rect 23792 6554 23816 6556
rect 23872 6554 23896 6556
rect 23952 6554 23976 6556
rect 23712 6502 23722 6554
rect 23966 6502 23976 6554
rect 23712 6500 23736 6502
rect 23792 6500 23816 6502
rect 23872 6500 23896 6502
rect 23952 6500 23976 6502
rect 23656 6491 24032 6500
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23572 6452 23624 6458
rect 24136 6440 24164 8366
rect 24676 7812 24728 7818
rect 24676 7754 24728 7760
rect 24688 7342 24716 7754
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 23572 6394 23624 6400
rect 23952 6412 24164 6440
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22916 6012 23292 6021
rect 22972 6010 22996 6012
rect 23052 6010 23076 6012
rect 23132 6010 23156 6012
rect 23212 6010 23236 6012
rect 22972 5958 22982 6010
rect 23226 5958 23236 6010
rect 22972 5956 22996 5958
rect 23052 5956 23076 5958
rect 23132 5956 23156 5958
rect 23212 5956 23236 5958
rect 22916 5947 23292 5956
rect 23584 5914 23612 6394
rect 23952 6254 23980 6412
rect 24032 6316 24084 6322
rect 24228 6304 24256 6734
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24084 6276 24256 6304
rect 24032 6258 24084 6264
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23656 5468 24032 5477
rect 23712 5466 23736 5468
rect 23792 5466 23816 5468
rect 23872 5466 23896 5468
rect 23952 5466 23976 5468
rect 23712 5414 23722 5466
rect 23966 5414 23976 5466
rect 23712 5412 23736 5414
rect 23792 5412 23816 5414
rect 23872 5412 23896 5414
rect 23952 5412 23976 5414
rect 23656 5403 24032 5412
rect 22916 4924 23292 4933
rect 22972 4922 22996 4924
rect 23052 4922 23076 4924
rect 23132 4922 23156 4924
rect 23212 4922 23236 4924
rect 22972 4870 22982 4922
rect 23226 4870 23236 4922
rect 22972 4868 22996 4870
rect 23052 4868 23076 4870
rect 23132 4868 23156 4870
rect 23212 4868 23236 4870
rect 22916 4859 23292 4868
rect 24228 4554 24256 6276
rect 24320 5710 24348 6326
rect 24596 6322 24624 6734
rect 24872 6458 24900 7346
rect 24964 6866 24992 8842
rect 25148 8566 25176 9046
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25148 7342 25176 7482
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24780 6186 24808 6258
rect 24872 6254 24900 6394
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24780 5914 24808 6122
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24768 5908 24820 5914
rect 24768 5850 24820 5856
rect 24780 5710 24808 5850
rect 24872 5778 24900 6054
rect 25148 5778 25176 7278
rect 25240 7002 25268 9522
rect 25424 7546 25452 10542
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25700 9586 25728 9998
rect 25792 9586 25820 12038
rect 26068 11354 26096 17070
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26160 15570 26188 16050
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 26160 12918 26188 13670
rect 26252 13394 26280 15846
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26344 14006 26372 15302
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26436 14414 26464 14758
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 26068 10810 26096 11290
rect 26056 10804 26108 10810
rect 26056 10746 26108 10752
rect 26148 10056 26200 10062
rect 26148 9998 26200 10004
rect 26160 9625 26188 9998
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26344 9654 26372 9862
rect 26332 9648 26384 9654
rect 26146 9616 26202 9625
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25780 9580 25832 9586
rect 26332 9590 26384 9596
rect 26146 9551 26202 9560
rect 25780 9522 25832 9528
rect 25596 9376 25648 9382
rect 25596 9318 25648 9324
rect 25608 8974 25636 9318
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25228 6996 25280 7002
rect 25228 6938 25280 6944
rect 25700 6866 25728 9522
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 25792 9042 25820 9318
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25792 7818 25820 8774
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 25780 7812 25832 7818
rect 25780 7754 25832 7760
rect 25688 6860 25740 6866
rect 25688 6802 25740 6808
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 25240 5710 25268 6326
rect 25332 6118 25360 6734
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25424 6361 25452 6394
rect 25410 6352 25466 6361
rect 25410 6287 25466 6296
rect 25516 6186 25544 6598
rect 25608 6390 25636 6598
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25504 6180 25556 6186
rect 25504 6122 25556 6128
rect 25608 6118 25636 6326
rect 25700 6322 25728 6666
rect 25976 6361 26004 7890
rect 26514 7576 26570 7585
rect 26514 7511 26516 7520
rect 26568 7511 26570 7520
rect 26516 7482 26568 7488
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26344 7313 26372 7346
rect 26330 7304 26386 7313
rect 26330 7239 26386 7248
rect 25962 6352 26018 6361
rect 25688 6316 25740 6322
rect 25962 6287 25964 6296
rect 25688 6258 25740 6264
rect 26016 6287 26018 6296
rect 25964 6258 26016 6264
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 25596 6112 25648 6118
rect 25596 6054 25648 6060
rect 25608 5846 25636 6054
rect 25596 5840 25648 5846
rect 25596 5782 25648 5788
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25596 5704 25648 5710
rect 25700 5692 25728 6258
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 26068 5846 26096 6054
rect 26056 5840 26108 5846
rect 26056 5782 26108 5788
rect 25648 5664 25728 5692
rect 25596 5646 25648 5652
rect 24216 4548 24268 4554
rect 24216 4490 24268 4496
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 22916 3836 23292 3845
rect 22972 3834 22996 3836
rect 23052 3834 23076 3836
rect 23132 3834 23156 3836
rect 23212 3834 23236 3836
rect 22972 3782 22982 3834
rect 23226 3782 23236 3834
rect 22972 3780 22996 3782
rect 23052 3780 23076 3782
rect 23132 3780 23156 3782
rect 23212 3780 23236 3782
rect 22916 3771 23292 3780
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22756 3398 22784 3538
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 23032 3058 23060 3470
rect 23492 3126 23520 4422
rect 23656 4380 24032 4389
rect 23712 4378 23736 4380
rect 23792 4378 23816 4380
rect 23872 4378 23896 4380
rect 23952 4378 23976 4380
rect 23712 4326 23722 4378
rect 23966 4326 23976 4378
rect 23712 4324 23736 4326
rect 23792 4324 23816 4326
rect 23872 4324 23896 4326
rect 23952 4324 23976 4326
rect 23656 4315 24032 4324
rect 24228 4214 24256 4490
rect 24216 4208 24268 4214
rect 24216 4150 24268 4156
rect 23656 3292 24032 3301
rect 23712 3290 23736 3292
rect 23792 3290 23816 3292
rect 23872 3290 23896 3292
rect 23952 3290 23976 3292
rect 23712 3238 23722 3290
rect 23966 3238 23976 3290
rect 23712 3236 23736 3238
rect 23792 3236 23816 3238
rect 23872 3236 23896 3238
rect 23952 3236 23976 3238
rect 23656 3227 24032 3236
rect 24320 3194 24348 5646
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 24412 4622 24440 5510
rect 25240 4622 25268 5510
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24412 4214 24440 4422
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 24952 4208 25004 4214
rect 24952 4150 25004 4156
rect 24964 3738 24992 4150
rect 25700 4146 25728 5664
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24308 3188 24360 3194
rect 24308 3130 24360 3136
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 24504 3058 24532 3334
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 22916 2748 23292 2757
rect 22972 2746 22996 2748
rect 23052 2746 23076 2748
rect 23132 2746 23156 2748
rect 23212 2746 23236 2748
rect 22972 2694 22982 2746
rect 23226 2694 23236 2746
rect 22972 2692 22996 2694
rect 23052 2692 23076 2694
rect 23132 2692 23156 2694
rect 23212 2692 23236 2694
rect 22916 2683 23292 2692
rect 19656 2204 20032 2213
rect 19712 2202 19736 2204
rect 19792 2202 19816 2204
rect 19872 2202 19896 2204
rect 19952 2202 19976 2204
rect 19712 2150 19722 2202
rect 19966 2150 19976 2202
rect 19712 2148 19736 2150
rect 19792 2148 19816 2150
rect 19872 2148 19896 2150
rect 19952 2148 19976 2150
rect 19656 2139 20032 2148
rect 23656 2204 24032 2213
rect 23712 2202 23736 2204
rect 23792 2202 23816 2204
rect 23872 2202 23896 2204
rect 23952 2202 23976 2204
rect 23712 2150 23722 2202
rect 23966 2150 23976 2202
rect 23712 2148 23736 2150
rect 23792 2148 23816 2150
rect 23872 2148 23896 2150
rect 23952 2148 23976 2150
rect 23656 2139 24032 2148
rect 5814 0 5870 800
rect 8390 0 8446 800
rect 12898 0 12954 800
rect 16118 0 16174 800
rect 19338 0 19394 800
<< via2 >>
rect 2916 27770 2972 27772
rect 2996 27770 3052 27772
rect 3076 27770 3132 27772
rect 3156 27770 3212 27772
rect 3236 27770 3292 27772
rect 2916 27718 2918 27770
rect 2918 27718 2970 27770
rect 2970 27718 2972 27770
rect 2996 27718 3034 27770
rect 3034 27718 3046 27770
rect 3046 27718 3052 27770
rect 3076 27718 3098 27770
rect 3098 27718 3110 27770
rect 3110 27718 3132 27770
rect 3156 27718 3162 27770
rect 3162 27718 3174 27770
rect 3174 27718 3212 27770
rect 3236 27718 3238 27770
rect 3238 27718 3290 27770
rect 3290 27718 3292 27770
rect 2916 27716 2972 27718
rect 2996 27716 3052 27718
rect 3076 27716 3132 27718
rect 3156 27716 3212 27718
rect 3236 27716 3292 27718
rect 6916 27770 6972 27772
rect 6996 27770 7052 27772
rect 7076 27770 7132 27772
rect 7156 27770 7212 27772
rect 7236 27770 7292 27772
rect 6916 27718 6918 27770
rect 6918 27718 6970 27770
rect 6970 27718 6972 27770
rect 6996 27718 7034 27770
rect 7034 27718 7046 27770
rect 7046 27718 7052 27770
rect 7076 27718 7098 27770
rect 7098 27718 7110 27770
rect 7110 27718 7132 27770
rect 7156 27718 7162 27770
rect 7162 27718 7174 27770
rect 7174 27718 7212 27770
rect 7236 27718 7238 27770
rect 7238 27718 7290 27770
rect 7290 27718 7292 27770
rect 6916 27716 6972 27718
rect 6996 27716 7052 27718
rect 7076 27716 7132 27718
rect 7156 27716 7212 27718
rect 7236 27716 7292 27718
rect 10916 27770 10972 27772
rect 10996 27770 11052 27772
rect 11076 27770 11132 27772
rect 11156 27770 11212 27772
rect 11236 27770 11292 27772
rect 10916 27718 10918 27770
rect 10918 27718 10970 27770
rect 10970 27718 10972 27770
rect 10996 27718 11034 27770
rect 11034 27718 11046 27770
rect 11046 27718 11052 27770
rect 11076 27718 11098 27770
rect 11098 27718 11110 27770
rect 11110 27718 11132 27770
rect 11156 27718 11162 27770
rect 11162 27718 11174 27770
rect 11174 27718 11212 27770
rect 11236 27718 11238 27770
rect 11238 27718 11290 27770
rect 11290 27718 11292 27770
rect 10916 27716 10972 27718
rect 10996 27716 11052 27718
rect 11076 27716 11132 27718
rect 11156 27716 11212 27718
rect 11236 27716 11292 27718
rect 14916 27770 14972 27772
rect 14996 27770 15052 27772
rect 15076 27770 15132 27772
rect 15156 27770 15212 27772
rect 15236 27770 15292 27772
rect 14916 27718 14918 27770
rect 14918 27718 14970 27770
rect 14970 27718 14972 27770
rect 14996 27718 15034 27770
rect 15034 27718 15046 27770
rect 15046 27718 15052 27770
rect 15076 27718 15098 27770
rect 15098 27718 15110 27770
rect 15110 27718 15132 27770
rect 15156 27718 15162 27770
rect 15162 27718 15174 27770
rect 15174 27718 15212 27770
rect 15236 27718 15238 27770
rect 15238 27718 15290 27770
rect 15290 27718 15292 27770
rect 14916 27716 14972 27718
rect 14996 27716 15052 27718
rect 15076 27716 15132 27718
rect 15156 27716 15212 27718
rect 15236 27716 15292 27718
rect 18916 27770 18972 27772
rect 18996 27770 19052 27772
rect 19076 27770 19132 27772
rect 19156 27770 19212 27772
rect 19236 27770 19292 27772
rect 18916 27718 18918 27770
rect 18918 27718 18970 27770
rect 18970 27718 18972 27770
rect 18996 27718 19034 27770
rect 19034 27718 19046 27770
rect 19046 27718 19052 27770
rect 19076 27718 19098 27770
rect 19098 27718 19110 27770
rect 19110 27718 19132 27770
rect 19156 27718 19162 27770
rect 19162 27718 19174 27770
rect 19174 27718 19212 27770
rect 19236 27718 19238 27770
rect 19238 27718 19290 27770
rect 19290 27718 19292 27770
rect 18916 27716 18972 27718
rect 18996 27716 19052 27718
rect 19076 27716 19132 27718
rect 19156 27716 19212 27718
rect 19236 27716 19292 27718
rect 3656 27226 3712 27228
rect 3736 27226 3792 27228
rect 3816 27226 3872 27228
rect 3896 27226 3952 27228
rect 3976 27226 4032 27228
rect 3656 27174 3658 27226
rect 3658 27174 3710 27226
rect 3710 27174 3712 27226
rect 3736 27174 3774 27226
rect 3774 27174 3786 27226
rect 3786 27174 3792 27226
rect 3816 27174 3838 27226
rect 3838 27174 3850 27226
rect 3850 27174 3872 27226
rect 3896 27174 3902 27226
rect 3902 27174 3914 27226
rect 3914 27174 3952 27226
rect 3976 27174 3978 27226
rect 3978 27174 4030 27226
rect 4030 27174 4032 27226
rect 3656 27172 3712 27174
rect 3736 27172 3792 27174
rect 3816 27172 3872 27174
rect 3896 27172 3952 27174
rect 3976 27172 4032 27174
rect 7656 27226 7712 27228
rect 7736 27226 7792 27228
rect 7816 27226 7872 27228
rect 7896 27226 7952 27228
rect 7976 27226 8032 27228
rect 7656 27174 7658 27226
rect 7658 27174 7710 27226
rect 7710 27174 7712 27226
rect 7736 27174 7774 27226
rect 7774 27174 7786 27226
rect 7786 27174 7792 27226
rect 7816 27174 7838 27226
rect 7838 27174 7850 27226
rect 7850 27174 7872 27226
rect 7896 27174 7902 27226
rect 7902 27174 7914 27226
rect 7914 27174 7952 27226
rect 7976 27174 7978 27226
rect 7978 27174 8030 27226
rect 8030 27174 8032 27226
rect 7656 27172 7712 27174
rect 7736 27172 7792 27174
rect 7816 27172 7872 27174
rect 7896 27172 7952 27174
rect 7976 27172 8032 27174
rect 2916 26682 2972 26684
rect 2996 26682 3052 26684
rect 3076 26682 3132 26684
rect 3156 26682 3212 26684
rect 3236 26682 3292 26684
rect 2916 26630 2918 26682
rect 2918 26630 2970 26682
rect 2970 26630 2972 26682
rect 2996 26630 3034 26682
rect 3034 26630 3046 26682
rect 3046 26630 3052 26682
rect 3076 26630 3098 26682
rect 3098 26630 3110 26682
rect 3110 26630 3132 26682
rect 3156 26630 3162 26682
rect 3162 26630 3174 26682
rect 3174 26630 3212 26682
rect 3236 26630 3238 26682
rect 3238 26630 3290 26682
rect 3290 26630 3292 26682
rect 2916 26628 2972 26630
rect 2996 26628 3052 26630
rect 3076 26628 3132 26630
rect 3156 26628 3212 26630
rect 3236 26628 3292 26630
rect 3422 26424 3478 26480
rect 2916 25594 2972 25596
rect 2996 25594 3052 25596
rect 3076 25594 3132 25596
rect 3156 25594 3212 25596
rect 3236 25594 3292 25596
rect 2916 25542 2918 25594
rect 2918 25542 2970 25594
rect 2970 25542 2972 25594
rect 2996 25542 3034 25594
rect 3034 25542 3046 25594
rect 3046 25542 3052 25594
rect 3076 25542 3098 25594
rect 3098 25542 3110 25594
rect 3110 25542 3132 25594
rect 3156 25542 3162 25594
rect 3162 25542 3174 25594
rect 3174 25542 3212 25594
rect 3236 25542 3238 25594
rect 3238 25542 3290 25594
rect 3290 25542 3292 25594
rect 2916 25540 2972 25542
rect 2996 25540 3052 25542
rect 3076 25540 3132 25542
rect 3156 25540 3212 25542
rect 3236 25540 3292 25542
rect 2916 24506 2972 24508
rect 2996 24506 3052 24508
rect 3076 24506 3132 24508
rect 3156 24506 3212 24508
rect 3236 24506 3292 24508
rect 2916 24454 2918 24506
rect 2918 24454 2970 24506
rect 2970 24454 2972 24506
rect 2996 24454 3034 24506
rect 3034 24454 3046 24506
rect 3046 24454 3052 24506
rect 3076 24454 3098 24506
rect 3098 24454 3110 24506
rect 3110 24454 3132 24506
rect 3156 24454 3162 24506
rect 3162 24454 3174 24506
rect 3174 24454 3212 24506
rect 3236 24454 3238 24506
rect 3238 24454 3290 24506
rect 3290 24454 3292 24506
rect 2916 24452 2972 24454
rect 2996 24452 3052 24454
rect 3076 24452 3132 24454
rect 3156 24452 3212 24454
rect 3236 24452 3292 24454
rect 2916 23418 2972 23420
rect 2996 23418 3052 23420
rect 3076 23418 3132 23420
rect 3156 23418 3212 23420
rect 3236 23418 3292 23420
rect 2916 23366 2918 23418
rect 2918 23366 2970 23418
rect 2970 23366 2972 23418
rect 2996 23366 3034 23418
rect 3034 23366 3046 23418
rect 3046 23366 3052 23418
rect 3076 23366 3098 23418
rect 3098 23366 3110 23418
rect 3110 23366 3132 23418
rect 3156 23366 3162 23418
rect 3162 23366 3174 23418
rect 3174 23366 3212 23418
rect 3236 23366 3238 23418
rect 3238 23366 3290 23418
rect 3290 23366 3292 23418
rect 2916 23364 2972 23366
rect 2996 23364 3052 23366
rect 3076 23364 3132 23366
rect 3156 23364 3212 23366
rect 3236 23364 3292 23366
rect 2916 22330 2972 22332
rect 2996 22330 3052 22332
rect 3076 22330 3132 22332
rect 3156 22330 3212 22332
rect 3236 22330 3292 22332
rect 2916 22278 2918 22330
rect 2918 22278 2970 22330
rect 2970 22278 2972 22330
rect 2996 22278 3034 22330
rect 3034 22278 3046 22330
rect 3046 22278 3052 22330
rect 3076 22278 3098 22330
rect 3098 22278 3110 22330
rect 3110 22278 3132 22330
rect 3156 22278 3162 22330
rect 3162 22278 3174 22330
rect 3174 22278 3212 22330
rect 3236 22278 3238 22330
rect 3238 22278 3290 22330
rect 3290 22278 3292 22330
rect 2916 22276 2972 22278
rect 2996 22276 3052 22278
rect 3076 22276 3132 22278
rect 3156 22276 3212 22278
rect 3236 22276 3292 22278
rect 2916 21242 2972 21244
rect 2996 21242 3052 21244
rect 3076 21242 3132 21244
rect 3156 21242 3212 21244
rect 3236 21242 3292 21244
rect 2916 21190 2918 21242
rect 2918 21190 2970 21242
rect 2970 21190 2972 21242
rect 2996 21190 3034 21242
rect 3034 21190 3046 21242
rect 3046 21190 3052 21242
rect 3076 21190 3098 21242
rect 3098 21190 3110 21242
rect 3110 21190 3132 21242
rect 3156 21190 3162 21242
rect 3162 21190 3174 21242
rect 3174 21190 3212 21242
rect 3236 21190 3238 21242
rect 3238 21190 3290 21242
rect 3290 21190 3292 21242
rect 2916 21188 2972 21190
rect 2996 21188 3052 21190
rect 3076 21188 3132 21190
rect 3156 21188 3212 21190
rect 3236 21188 3292 21190
rect 2916 20154 2972 20156
rect 2996 20154 3052 20156
rect 3076 20154 3132 20156
rect 3156 20154 3212 20156
rect 3236 20154 3292 20156
rect 2916 20102 2918 20154
rect 2918 20102 2970 20154
rect 2970 20102 2972 20154
rect 2996 20102 3034 20154
rect 3034 20102 3046 20154
rect 3046 20102 3052 20154
rect 3076 20102 3098 20154
rect 3098 20102 3110 20154
rect 3110 20102 3132 20154
rect 3156 20102 3162 20154
rect 3162 20102 3174 20154
rect 3174 20102 3212 20154
rect 3236 20102 3238 20154
rect 3238 20102 3290 20154
rect 3290 20102 3292 20154
rect 2916 20100 2972 20102
rect 2996 20100 3052 20102
rect 3076 20100 3132 20102
rect 3156 20100 3212 20102
rect 3236 20100 3292 20102
rect 1398 17720 1454 17776
rect 2916 19066 2972 19068
rect 2996 19066 3052 19068
rect 3076 19066 3132 19068
rect 3156 19066 3212 19068
rect 3236 19066 3292 19068
rect 2916 19014 2918 19066
rect 2918 19014 2970 19066
rect 2970 19014 2972 19066
rect 2996 19014 3034 19066
rect 3034 19014 3046 19066
rect 3046 19014 3052 19066
rect 3076 19014 3098 19066
rect 3098 19014 3110 19066
rect 3110 19014 3132 19066
rect 3156 19014 3162 19066
rect 3162 19014 3174 19066
rect 3174 19014 3212 19066
rect 3236 19014 3238 19066
rect 3238 19014 3290 19066
rect 3290 19014 3292 19066
rect 2916 19012 2972 19014
rect 2996 19012 3052 19014
rect 3076 19012 3132 19014
rect 3156 19012 3212 19014
rect 3236 19012 3292 19014
rect 2916 17978 2972 17980
rect 2996 17978 3052 17980
rect 3076 17978 3132 17980
rect 3156 17978 3212 17980
rect 3236 17978 3292 17980
rect 2916 17926 2918 17978
rect 2918 17926 2970 17978
rect 2970 17926 2972 17978
rect 2996 17926 3034 17978
rect 3034 17926 3046 17978
rect 3046 17926 3052 17978
rect 3076 17926 3098 17978
rect 3098 17926 3110 17978
rect 3110 17926 3132 17978
rect 3156 17926 3162 17978
rect 3162 17926 3174 17978
rect 3174 17926 3212 17978
rect 3236 17926 3238 17978
rect 3238 17926 3290 17978
rect 3290 17926 3292 17978
rect 2916 17924 2972 17926
rect 2996 17924 3052 17926
rect 3076 17924 3132 17926
rect 3156 17924 3212 17926
rect 3236 17924 3292 17926
rect 2916 16890 2972 16892
rect 2996 16890 3052 16892
rect 3076 16890 3132 16892
rect 3156 16890 3212 16892
rect 3236 16890 3292 16892
rect 2916 16838 2918 16890
rect 2918 16838 2970 16890
rect 2970 16838 2972 16890
rect 2996 16838 3034 16890
rect 3034 16838 3046 16890
rect 3046 16838 3052 16890
rect 3076 16838 3098 16890
rect 3098 16838 3110 16890
rect 3110 16838 3132 16890
rect 3156 16838 3162 16890
rect 3162 16838 3174 16890
rect 3174 16838 3212 16890
rect 3236 16838 3238 16890
rect 3238 16838 3290 16890
rect 3290 16838 3292 16890
rect 2916 16836 2972 16838
rect 2996 16836 3052 16838
rect 3076 16836 3132 16838
rect 3156 16836 3212 16838
rect 3236 16836 3292 16838
rect 2916 15802 2972 15804
rect 2996 15802 3052 15804
rect 3076 15802 3132 15804
rect 3156 15802 3212 15804
rect 3236 15802 3292 15804
rect 2916 15750 2918 15802
rect 2918 15750 2970 15802
rect 2970 15750 2972 15802
rect 2996 15750 3034 15802
rect 3034 15750 3046 15802
rect 3046 15750 3052 15802
rect 3076 15750 3098 15802
rect 3098 15750 3110 15802
rect 3110 15750 3132 15802
rect 3156 15750 3162 15802
rect 3162 15750 3174 15802
rect 3174 15750 3212 15802
rect 3236 15750 3238 15802
rect 3238 15750 3290 15802
rect 3290 15750 3292 15802
rect 2916 15748 2972 15750
rect 2996 15748 3052 15750
rect 3076 15748 3132 15750
rect 3156 15748 3212 15750
rect 3236 15748 3292 15750
rect 3656 26138 3712 26140
rect 3736 26138 3792 26140
rect 3816 26138 3872 26140
rect 3896 26138 3952 26140
rect 3976 26138 4032 26140
rect 3656 26086 3658 26138
rect 3658 26086 3710 26138
rect 3710 26086 3712 26138
rect 3736 26086 3774 26138
rect 3774 26086 3786 26138
rect 3786 26086 3792 26138
rect 3816 26086 3838 26138
rect 3838 26086 3850 26138
rect 3850 26086 3872 26138
rect 3896 26086 3902 26138
rect 3902 26086 3914 26138
rect 3914 26086 3952 26138
rect 3976 26086 3978 26138
rect 3978 26086 4030 26138
rect 4030 26086 4032 26138
rect 3656 26084 3712 26086
rect 3736 26084 3792 26086
rect 3816 26084 3872 26086
rect 3896 26084 3952 26086
rect 3976 26084 4032 26086
rect 6916 26682 6972 26684
rect 6996 26682 7052 26684
rect 7076 26682 7132 26684
rect 7156 26682 7212 26684
rect 7236 26682 7292 26684
rect 6916 26630 6918 26682
rect 6918 26630 6970 26682
rect 6970 26630 6972 26682
rect 6996 26630 7034 26682
rect 7034 26630 7046 26682
rect 7046 26630 7052 26682
rect 7076 26630 7098 26682
rect 7098 26630 7110 26682
rect 7110 26630 7132 26682
rect 7156 26630 7162 26682
rect 7162 26630 7174 26682
rect 7174 26630 7212 26682
rect 7236 26630 7238 26682
rect 7238 26630 7290 26682
rect 7290 26630 7292 26682
rect 6916 26628 6972 26630
rect 6996 26628 7052 26630
rect 7076 26628 7132 26630
rect 7156 26628 7212 26630
rect 7236 26628 7292 26630
rect 3656 25050 3712 25052
rect 3736 25050 3792 25052
rect 3816 25050 3872 25052
rect 3896 25050 3952 25052
rect 3976 25050 4032 25052
rect 3656 24998 3658 25050
rect 3658 24998 3710 25050
rect 3710 24998 3712 25050
rect 3736 24998 3774 25050
rect 3774 24998 3786 25050
rect 3786 24998 3792 25050
rect 3816 24998 3838 25050
rect 3838 24998 3850 25050
rect 3850 24998 3872 25050
rect 3896 24998 3902 25050
rect 3902 24998 3914 25050
rect 3914 24998 3952 25050
rect 3976 24998 3978 25050
rect 3978 24998 4030 25050
rect 4030 24998 4032 25050
rect 3656 24996 3712 24998
rect 3736 24996 3792 24998
rect 3816 24996 3872 24998
rect 3896 24996 3952 24998
rect 3976 24996 4032 24998
rect 3656 23962 3712 23964
rect 3736 23962 3792 23964
rect 3816 23962 3872 23964
rect 3896 23962 3952 23964
rect 3976 23962 4032 23964
rect 3656 23910 3658 23962
rect 3658 23910 3710 23962
rect 3710 23910 3712 23962
rect 3736 23910 3774 23962
rect 3774 23910 3786 23962
rect 3786 23910 3792 23962
rect 3816 23910 3838 23962
rect 3838 23910 3850 23962
rect 3850 23910 3872 23962
rect 3896 23910 3902 23962
rect 3902 23910 3914 23962
rect 3914 23910 3952 23962
rect 3976 23910 3978 23962
rect 3978 23910 4030 23962
rect 4030 23910 4032 23962
rect 3656 23908 3712 23910
rect 3736 23908 3792 23910
rect 3816 23908 3872 23910
rect 3896 23908 3952 23910
rect 3976 23908 4032 23910
rect 3656 22874 3712 22876
rect 3736 22874 3792 22876
rect 3816 22874 3872 22876
rect 3896 22874 3952 22876
rect 3976 22874 4032 22876
rect 3656 22822 3658 22874
rect 3658 22822 3710 22874
rect 3710 22822 3712 22874
rect 3736 22822 3774 22874
rect 3774 22822 3786 22874
rect 3786 22822 3792 22874
rect 3816 22822 3838 22874
rect 3838 22822 3850 22874
rect 3850 22822 3872 22874
rect 3896 22822 3902 22874
rect 3902 22822 3914 22874
rect 3914 22822 3952 22874
rect 3976 22822 3978 22874
rect 3978 22822 4030 22874
rect 4030 22822 4032 22874
rect 3656 22820 3712 22822
rect 3736 22820 3792 22822
rect 3816 22820 3872 22822
rect 3896 22820 3952 22822
rect 3976 22820 4032 22822
rect 3656 21786 3712 21788
rect 3736 21786 3792 21788
rect 3816 21786 3872 21788
rect 3896 21786 3952 21788
rect 3976 21786 4032 21788
rect 3656 21734 3658 21786
rect 3658 21734 3710 21786
rect 3710 21734 3712 21786
rect 3736 21734 3774 21786
rect 3774 21734 3786 21786
rect 3786 21734 3792 21786
rect 3816 21734 3838 21786
rect 3838 21734 3850 21786
rect 3850 21734 3872 21786
rect 3896 21734 3902 21786
rect 3902 21734 3914 21786
rect 3914 21734 3952 21786
rect 3976 21734 3978 21786
rect 3978 21734 4030 21786
rect 4030 21734 4032 21786
rect 3656 21732 3712 21734
rect 3736 21732 3792 21734
rect 3816 21732 3872 21734
rect 3896 21732 3952 21734
rect 3976 21732 4032 21734
rect 3656 20698 3712 20700
rect 3736 20698 3792 20700
rect 3816 20698 3872 20700
rect 3896 20698 3952 20700
rect 3976 20698 4032 20700
rect 3656 20646 3658 20698
rect 3658 20646 3710 20698
rect 3710 20646 3712 20698
rect 3736 20646 3774 20698
rect 3774 20646 3786 20698
rect 3786 20646 3792 20698
rect 3816 20646 3838 20698
rect 3838 20646 3850 20698
rect 3850 20646 3872 20698
rect 3896 20646 3902 20698
rect 3902 20646 3914 20698
rect 3914 20646 3952 20698
rect 3976 20646 3978 20698
rect 3978 20646 4030 20698
rect 4030 20646 4032 20698
rect 3656 20644 3712 20646
rect 3736 20644 3792 20646
rect 3816 20644 3872 20646
rect 3896 20644 3952 20646
rect 3976 20644 4032 20646
rect 3656 19610 3712 19612
rect 3736 19610 3792 19612
rect 3816 19610 3872 19612
rect 3896 19610 3952 19612
rect 3976 19610 4032 19612
rect 3656 19558 3658 19610
rect 3658 19558 3710 19610
rect 3710 19558 3712 19610
rect 3736 19558 3774 19610
rect 3774 19558 3786 19610
rect 3786 19558 3792 19610
rect 3816 19558 3838 19610
rect 3838 19558 3850 19610
rect 3850 19558 3872 19610
rect 3896 19558 3902 19610
rect 3902 19558 3914 19610
rect 3914 19558 3952 19610
rect 3976 19558 3978 19610
rect 3978 19558 4030 19610
rect 4030 19558 4032 19610
rect 3656 19556 3712 19558
rect 3736 19556 3792 19558
rect 3816 19556 3872 19558
rect 3896 19556 3952 19558
rect 3976 19556 4032 19558
rect 3656 18522 3712 18524
rect 3736 18522 3792 18524
rect 3816 18522 3872 18524
rect 3896 18522 3952 18524
rect 3976 18522 4032 18524
rect 3656 18470 3658 18522
rect 3658 18470 3710 18522
rect 3710 18470 3712 18522
rect 3736 18470 3774 18522
rect 3774 18470 3786 18522
rect 3786 18470 3792 18522
rect 3816 18470 3838 18522
rect 3838 18470 3850 18522
rect 3850 18470 3872 18522
rect 3896 18470 3902 18522
rect 3902 18470 3914 18522
rect 3914 18470 3952 18522
rect 3976 18470 3978 18522
rect 3978 18470 4030 18522
rect 4030 18470 4032 18522
rect 3656 18468 3712 18470
rect 3736 18468 3792 18470
rect 3816 18468 3872 18470
rect 3896 18468 3952 18470
rect 3976 18468 4032 18470
rect 3656 17434 3712 17436
rect 3736 17434 3792 17436
rect 3816 17434 3872 17436
rect 3896 17434 3952 17436
rect 3976 17434 4032 17436
rect 3656 17382 3658 17434
rect 3658 17382 3710 17434
rect 3710 17382 3712 17434
rect 3736 17382 3774 17434
rect 3774 17382 3786 17434
rect 3786 17382 3792 17434
rect 3816 17382 3838 17434
rect 3838 17382 3850 17434
rect 3850 17382 3872 17434
rect 3896 17382 3902 17434
rect 3902 17382 3914 17434
rect 3914 17382 3952 17434
rect 3976 17382 3978 17434
rect 3978 17382 4030 17434
rect 4030 17382 4032 17434
rect 3656 17380 3712 17382
rect 3736 17380 3792 17382
rect 3816 17380 3872 17382
rect 3896 17380 3952 17382
rect 3976 17380 4032 17382
rect 2916 14714 2972 14716
rect 2996 14714 3052 14716
rect 3076 14714 3132 14716
rect 3156 14714 3212 14716
rect 3236 14714 3292 14716
rect 2916 14662 2918 14714
rect 2918 14662 2970 14714
rect 2970 14662 2972 14714
rect 2996 14662 3034 14714
rect 3034 14662 3046 14714
rect 3046 14662 3052 14714
rect 3076 14662 3098 14714
rect 3098 14662 3110 14714
rect 3110 14662 3132 14714
rect 3156 14662 3162 14714
rect 3162 14662 3174 14714
rect 3174 14662 3212 14714
rect 3236 14662 3238 14714
rect 3238 14662 3290 14714
rect 3290 14662 3292 14714
rect 2916 14660 2972 14662
rect 2996 14660 3052 14662
rect 3076 14660 3132 14662
rect 3156 14660 3212 14662
rect 3236 14660 3292 14662
rect 3422 15000 3478 15056
rect 2916 13626 2972 13628
rect 2996 13626 3052 13628
rect 3076 13626 3132 13628
rect 3156 13626 3212 13628
rect 3236 13626 3292 13628
rect 2916 13574 2918 13626
rect 2918 13574 2970 13626
rect 2970 13574 2972 13626
rect 2996 13574 3034 13626
rect 3034 13574 3046 13626
rect 3046 13574 3052 13626
rect 3076 13574 3098 13626
rect 3098 13574 3110 13626
rect 3110 13574 3132 13626
rect 3156 13574 3162 13626
rect 3162 13574 3174 13626
rect 3174 13574 3212 13626
rect 3236 13574 3238 13626
rect 3238 13574 3290 13626
rect 3290 13574 3292 13626
rect 2916 13572 2972 13574
rect 2996 13572 3052 13574
rect 3076 13572 3132 13574
rect 3156 13572 3212 13574
rect 3236 13572 3292 13574
rect 846 12844 902 12880
rect 846 12824 848 12844
rect 848 12824 900 12844
rect 900 12824 902 12844
rect 2916 12538 2972 12540
rect 2996 12538 3052 12540
rect 3076 12538 3132 12540
rect 3156 12538 3212 12540
rect 3236 12538 3292 12540
rect 2916 12486 2918 12538
rect 2918 12486 2970 12538
rect 2970 12486 2972 12538
rect 2996 12486 3034 12538
rect 3034 12486 3046 12538
rect 3046 12486 3052 12538
rect 3076 12486 3098 12538
rect 3098 12486 3110 12538
rect 3110 12486 3132 12538
rect 3156 12486 3162 12538
rect 3162 12486 3174 12538
rect 3174 12486 3212 12538
rect 3236 12486 3238 12538
rect 3238 12486 3290 12538
rect 3290 12486 3292 12538
rect 2916 12484 2972 12486
rect 2996 12484 3052 12486
rect 3076 12484 3132 12486
rect 3156 12484 3212 12486
rect 3236 12484 3292 12486
rect 2916 11450 2972 11452
rect 2996 11450 3052 11452
rect 3076 11450 3132 11452
rect 3156 11450 3212 11452
rect 3236 11450 3292 11452
rect 2916 11398 2918 11450
rect 2918 11398 2970 11450
rect 2970 11398 2972 11450
rect 2996 11398 3034 11450
rect 3034 11398 3046 11450
rect 3046 11398 3052 11450
rect 3076 11398 3098 11450
rect 3098 11398 3110 11450
rect 3110 11398 3132 11450
rect 3156 11398 3162 11450
rect 3162 11398 3174 11450
rect 3174 11398 3212 11450
rect 3236 11398 3238 11450
rect 3238 11398 3290 11450
rect 3290 11398 3292 11450
rect 2916 11396 2972 11398
rect 2996 11396 3052 11398
rect 3076 11396 3132 11398
rect 3156 11396 3212 11398
rect 3236 11396 3292 11398
rect 2916 10362 2972 10364
rect 2996 10362 3052 10364
rect 3076 10362 3132 10364
rect 3156 10362 3212 10364
rect 3236 10362 3292 10364
rect 2916 10310 2918 10362
rect 2918 10310 2970 10362
rect 2970 10310 2972 10362
rect 2996 10310 3034 10362
rect 3034 10310 3046 10362
rect 3046 10310 3052 10362
rect 3076 10310 3098 10362
rect 3098 10310 3110 10362
rect 3110 10310 3132 10362
rect 3156 10310 3162 10362
rect 3162 10310 3174 10362
rect 3174 10310 3212 10362
rect 3236 10310 3238 10362
rect 3238 10310 3290 10362
rect 3290 10310 3292 10362
rect 2916 10308 2972 10310
rect 2996 10308 3052 10310
rect 3076 10308 3132 10310
rect 3156 10308 3212 10310
rect 3236 10308 3292 10310
rect 2686 9968 2742 10024
rect 1398 9560 1454 9616
rect 2916 9274 2972 9276
rect 2996 9274 3052 9276
rect 3076 9274 3132 9276
rect 3156 9274 3212 9276
rect 3236 9274 3292 9276
rect 2916 9222 2918 9274
rect 2918 9222 2970 9274
rect 2970 9222 2972 9274
rect 2996 9222 3034 9274
rect 3034 9222 3046 9274
rect 3046 9222 3052 9274
rect 3076 9222 3098 9274
rect 3098 9222 3110 9274
rect 3110 9222 3132 9274
rect 3156 9222 3162 9274
rect 3162 9222 3174 9274
rect 3174 9222 3212 9274
rect 3236 9222 3238 9274
rect 3238 9222 3290 9274
rect 3290 9222 3292 9274
rect 2916 9220 2972 9222
rect 2996 9220 3052 9222
rect 3076 9220 3132 9222
rect 3156 9220 3212 9222
rect 3236 9220 3292 9222
rect 3656 16346 3712 16348
rect 3736 16346 3792 16348
rect 3816 16346 3872 16348
rect 3896 16346 3952 16348
rect 3976 16346 4032 16348
rect 3656 16294 3658 16346
rect 3658 16294 3710 16346
rect 3710 16294 3712 16346
rect 3736 16294 3774 16346
rect 3774 16294 3786 16346
rect 3786 16294 3792 16346
rect 3816 16294 3838 16346
rect 3838 16294 3850 16346
rect 3850 16294 3872 16346
rect 3896 16294 3902 16346
rect 3902 16294 3914 16346
rect 3914 16294 3952 16346
rect 3976 16294 3978 16346
rect 3978 16294 4030 16346
rect 4030 16294 4032 16346
rect 3656 16292 3712 16294
rect 3736 16292 3792 16294
rect 3816 16292 3872 16294
rect 3896 16292 3952 16294
rect 3976 16292 4032 16294
rect 3656 15258 3712 15260
rect 3736 15258 3792 15260
rect 3816 15258 3872 15260
rect 3896 15258 3952 15260
rect 3976 15258 4032 15260
rect 3656 15206 3658 15258
rect 3658 15206 3710 15258
rect 3710 15206 3712 15258
rect 3736 15206 3774 15258
rect 3774 15206 3786 15258
rect 3786 15206 3792 15258
rect 3816 15206 3838 15258
rect 3838 15206 3850 15258
rect 3850 15206 3872 15258
rect 3896 15206 3902 15258
rect 3902 15206 3914 15258
rect 3914 15206 3952 15258
rect 3976 15206 3978 15258
rect 3978 15206 4030 15258
rect 4030 15206 4032 15258
rect 3656 15204 3712 15206
rect 3736 15204 3792 15206
rect 3816 15204 3872 15206
rect 3896 15204 3952 15206
rect 3976 15204 4032 15206
rect 3656 14170 3712 14172
rect 3736 14170 3792 14172
rect 3816 14170 3872 14172
rect 3896 14170 3952 14172
rect 3976 14170 4032 14172
rect 3656 14118 3658 14170
rect 3658 14118 3710 14170
rect 3710 14118 3712 14170
rect 3736 14118 3774 14170
rect 3774 14118 3786 14170
rect 3786 14118 3792 14170
rect 3816 14118 3838 14170
rect 3838 14118 3850 14170
rect 3850 14118 3872 14170
rect 3896 14118 3902 14170
rect 3902 14118 3914 14170
rect 3914 14118 3952 14170
rect 3976 14118 3978 14170
rect 3978 14118 4030 14170
rect 4030 14118 4032 14170
rect 3656 14116 3712 14118
rect 3736 14116 3792 14118
rect 3816 14116 3872 14118
rect 3896 14116 3952 14118
rect 3976 14116 4032 14118
rect 3656 13082 3712 13084
rect 3736 13082 3792 13084
rect 3816 13082 3872 13084
rect 3896 13082 3952 13084
rect 3976 13082 4032 13084
rect 3656 13030 3658 13082
rect 3658 13030 3710 13082
rect 3710 13030 3712 13082
rect 3736 13030 3774 13082
rect 3774 13030 3786 13082
rect 3786 13030 3792 13082
rect 3816 13030 3838 13082
rect 3838 13030 3850 13082
rect 3850 13030 3872 13082
rect 3896 13030 3902 13082
rect 3902 13030 3914 13082
rect 3914 13030 3952 13082
rect 3976 13030 3978 13082
rect 3978 13030 4030 13082
rect 4030 13030 4032 13082
rect 3656 13028 3712 13030
rect 3736 13028 3792 13030
rect 3816 13028 3872 13030
rect 3896 13028 3952 13030
rect 3976 13028 4032 13030
rect 3656 11994 3712 11996
rect 3736 11994 3792 11996
rect 3816 11994 3872 11996
rect 3896 11994 3952 11996
rect 3976 11994 4032 11996
rect 3656 11942 3658 11994
rect 3658 11942 3710 11994
rect 3710 11942 3712 11994
rect 3736 11942 3774 11994
rect 3774 11942 3786 11994
rect 3786 11942 3792 11994
rect 3816 11942 3838 11994
rect 3838 11942 3850 11994
rect 3850 11942 3872 11994
rect 3896 11942 3902 11994
rect 3902 11942 3914 11994
rect 3914 11942 3952 11994
rect 3976 11942 3978 11994
rect 3978 11942 4030 11994
rect 4030 11942 4032 11994
rect 3656 11940 3712 11942
rect 3736 11940 3792 11942
rect 3816 11940 3872 11942
rect 3896 11940 3952 11942
rect 3976 11940 4032 11942
rect 3698 11636 3700 11656
rect 3700 11636 3752 11656
rect 3752 11636 3754 11656
rect 3698 11600 3754 11636
rect 3656 10906 3712 10908
rect 3736 10906 3792 10908
rect 3816 10906 3872 10908
rect 3896 10906 3952 10908
rect 3976 10906 4032 10908
rect 3656 10854 3658 10906
rect 3658 10854 3710 10906
rect 3710 10854 3712 10906
rect 3736 10854 3774 10906
rect 3774 10854 3786 10906
rect 3786 10854 3792 10906
rect 3816 10854 3838 10906
rect 3838 10854 3850 10906
rect 3850 10854 3872 10906
rect 3896 10854 3902 10906
rect 3902 10854 3914 10906
rect 3914 10854 3952 10906
rect 3976 10854 3978 10906
rect 3978 10854 4030 10906
rect 4030 10854 4032 10906
rect 3656 10852 3712 10854
rect 3736 10852 3792 10854
rect 3816 10852 3872 10854
rect 3896 10852 3952 10854
rect 3976 10852 4032 10854
rect 5354 22072 5410 22128
rect 5262 19352 5318 19408
rect 6916 25594 6972 25596
rect 6996 25594 7052 25596
rect 7076 25594 7132 25596
rect 7156 25594 7212 25596
rect 7236 25594 7292 25596
rect 6916 25542 6918 25594
rect 6918 25542 6970 25594
rect 6970 25542 6972 25594
rect 6996 25542 7034 25594
rect 7034 25542 7046 25594
rect 7046 25542 7052 25594
rect 7076 25542 7098 25594
rect 7098 25542 7110 25594
rect 7110 25542 7132 25594
rect 7156 25542 7162 25594
rect 7162 25542 7174 25594
rect 7174 25542 7212 25594
rect 7236 25542 7238 25594
rect 7238 25542 7290 25594
rect 7290 25542 7292 25594
rect 6916 25540 6972 25542
rect 6996 25540 7052 25542
rect 7076 25540 7132 25542
rect 7156 25540 7212 25542
rect 7236 25540 7292 25542
rect 7656 26138 7712 26140
rect 7736 26138 7792 26140
rect 7816 26138 7872 26140
rect 7896 26138 7952 26140
rect 7976 26138 8032 26140
rect 7656 26086 7658 26138
rect 7658 26086 7710 26138
rect 7710 26086 7712 26138
rect 7736 26086 7774 26138
rect 7774 26086 7786 26138
rect 7786 26086 7792 26138
rect 7816 26086 7838 26138
rect 7838 26086 7850 26138
rect 7850 26086 7872 26138
rect 7896 26086 7902 26138
rect 7902 26086 7914 26138
rect 7914 26086 7952 26138
rect 7976 26086 7978 26138
rect 7978 26086 8030 26138
rect 8030 26086 8032 26138
rect 7656 26084 7712 26086
rect 7736 26084 7792 26086
rect 7816 26084 7872 26086
rect 7896 26084 7952 26086
rect 7976 26084 8032 26086
rect 7656 25050 7712 25052
rect 7736 25050 7792 25052
rect 7816 25050 7872 25052
rect 7896 25050 7952 25052
rect 7976 25050 8032 25052
rect 7656 24998 7658 25050
rect 7658 24998 7710 25050
rect 7710 24998 7712 25050
rect 7736 24998 7774 25050
rect 7774 24998 7786 25050
rect 7786 24998 7792 25050
rect 7816 24998 7838 25050
rect 7838 24998 7850 25050
rect 7850 24998 7872 25050
rect 7896 24998 7902 25050
rect 7902 24998 7914 25050
rect 7914 24998 7952 25050
rect 7976 24998 7978 25050
rect 7978 24998 8030 25050
rect 8030 24998 8032 25050
rect 7656 24996 7712 24998
rect 7736 24996 7792 24998
rect 7816 24996 7872 24998
rect 7896 24996 7952 24998
rect 7976 24996 8032 24998
rect 6916 24506 6972 24508
rect 6996 24506 7052 24508
rect 7076 24506 7132 24508
rect 7156 24506 7212 24508
rect 7236 24506 7292 24508
rect 6916 24454 6918 24506
rect 6918 24454 6970 24506
rect 6970 24454 6972 24506
rect 6996 24454 7034 24506
rect 7034 24454 7046 24506
rect 7046 24454 7052 24506
rect 7076 24454 7098 24506
rect 7098 24454 7110 24506
rect 7110 24454 7132 24506
rect 7156 24454 7162 24506
rect 7162 24454 7174 24506
rect 7174 24454 7212 24506
rect 7236 24454 7238 24506
rect 7238 24454 7290 24506
rect 7290 24454 7292 24506
rect 6916 24452 6972 24454
rect 6996 24452 7052 24454
rect 7076 24452 7132 24454
rect 7156 24452 7212 24454
rect 7236 24452 7292 24454
rect 6916 23418 6972 23420
rect 6996 23418 7052 23420
rect 7076 23418 7132 23420
rect 7156 23418 7212 23420
rect 7236 23418 7292 23420
rect 6916 23366 6918 23418
rect 6918 23366 6970 23418
rect 6970 23366 6972 23418
rect 6996 23366 7034 23418
rect 7034 23366 7046 23418
rect 7046 23366 7052 23418
rect 7076 23366 7098 23418
rect 7098 23366 7110 23418
rect 7110 23366 7132 23418
rect 7156 23366 7162 23418
rect 7162 23366 7174 23418
rect 7174 23366 7212 23418
rect 7236 23366 7238 23418
rect 7238 23366 7290 23418
rect 7290 23366 7292 23418
rect 6916 23364 6972 23366
rect 6996 23364 7052 23366
rect 7076 23364 7132 23366
rect 7156 23364 7212 23366
rect 7236 23364 7292 23366
rect 7656 23962 7712 23964
rect 7736 23962 7792 23964
rect 7816 23962 7872 23964
rect 7896 23962 7952 23964
rect 7976 23962 8032 23964
rect 7656 23910 7658 23962
rect 7658 23910 7710 23962
rect 7710 23910 7712 23962
rect 7736 23910 7774 23962
rect 7774 23910 7786 23962
rect 7786 23910 7792 23962
rect 7816 23910 7838 23962
rect 7838 23910 7850 23962
rect 7850 23910 7872 23962
rect 7896 23910 7902 23962
rect 7902 23910 7914 23962
rect 7914 23910 7952 23962
rect 7976 23910 7978 23962
rect 7978 23910 8030 23962
rect 8030 23910 8032 23962
rect 7656 23908 7712 23910
rect 7736 23908 7792 23910
rect 7816 23908 7872 23910
rect 7896 23908 7952 23910
rect 7976 23908 8032 23910
rect 5446 19372 5502 19408
rect 5446 19352 5448 19372
rect 5448 19352 5500 19372
rect 5500 19352 5502 19372
rect 4710 12824 4766 12880
rect 5262 12824 5318 12880
rect 6916 22330 6972 22332
rect 6996 22330 7052 22332
rect 7076 22330 7132 22332
rect 7156 22330 7212 22332
rect 7236 22330 7292 22332
rect 6916 22278 6918 22330
rect 6918 22278 6970 22330
rect 6970 22278 6972 22330
rect 6996 22278 7034 22330
rect 7034 22278 7046 22330
rect 7046 22278 7052 22330
rect 7076 22278 7098 22330
rect 7098 22278 7110 22330
rect 7110 22278 7132 22330
rect 7156 22278 7162 22330
rect 7162 22278 7174 22330
rect 7174 22278 7212 22330
rect 7236 22278 7238 22330
rect 7238 22278 7290 22330
rect 7290 22278 7292 22330
rect 6916 22276 6972 22278
rect 6996 22276 7052 22278
rect 7076 22276 7132 22278
rect 7156 22276 7212 22278
rect 7236 22276 7292 22278
rect 5354 12416 5410 12472
rect 3514 9968 3570 10024
rect 3656 9818 3712 9820
rect 3736 9818 3792 9820
rect 3816 9818 3872 9820
rect 3896 9818 3952 9820
rect 3976 9818 4032 9820
rect 3656 9766 3658 9818
rect 3658 9766 3710 9818
rect 3710 9766 3712 9818
rect 3736 9766 3774 9818
rect 3774 9766 3786 9818
rect 3786 9766 3792 9818
rect 3816 9766 3838 9818
rect 3838 9766 3850 9818
rect 3850 9766 3872 9818
rect 3896 9766 3902 9818
rect 3902 9766 3914 9818
rect 3914 9766 3952 9818
rect 3976 9766 3978 9818
rect 3978 9766 4030 9818
rect 4030 9766 4032 9818
rect 3656 9764 3712 9766
rect 3736 9764 3792 9766
rect 3816 9764 3872 9766
rect 3896 9764 3952 9766
rect 3976 9764 4032 9766
rect 3656 8730 3712 8732
rect 3736 8730 3792 8732
rect 3816 8730 3872 8732
rect 3896 8730 3952 8732
rect 3976 8730 4032 8732
rect 3656 8678 3658 8730
rect 3658 8678 3710 8730
rect 3710 8678 3712 8730
rect 3736 8678 3774 8730
rect 3774 8678 3786 8730
rect 3786 8678 3792 8730
rect 3816 8678 3838 8730
rect 3838 8678 3850 8730
rect 3850 8678 3872 8730
rect 3896 8678 3902 8730
rect 3902 8678 3914 8730
rect 3914 8678 3952 8730
rect 3976 8678 3978 8730
rect 3978 8678 4030 8730
rect 4030 8678 4032 8730
rect 3656 8676 3712 8678
rect 3736 8676 3792 8678
rect 3816 8676 3872 8678
rect 3896 8676 3952 8678
rect 3976 8676 4032 8678
rect 2916 8186 2972 8188
rect 2996 8186 3052 8188
rect 3076 8186 3132 8188
rect 3156 8186 3212 8188
rect 3236 8186 3292 8188
rect 2916 8134 2918 8186
rect 2918 8134 2970 8186
rect 2970 8134 2972 8186
rect 2996 8134 3034 8186
rect 3034 8134 3046 8186
rect 3046 8134 3052 8186
rect 3076 8134 3098 8186
rect 3098 8134 3110 8186
rect 3110 8134 3132 8186
rect 3156 8134 3162 8186
rect 3162 8134 3174 8186
rect 3174 8134 3212 8186
rect 3236 8134 3238 8186
rect 3238 8134 3290 8186
rect 3290 8134 3292 8186
rect 2916 8132 2972 8134
rect 2996 8132 3052 8134
rect 3076 8132 3132 8134
rect 3156 8132 3212 8134
rect 3236 8132 3292 8134
rect 3656 7642 3712 7644
rect 3736 7642 3792 7644
rect 3816 7642 3872 7644
rect 3896 7642 3952 7644
rect 3976 7642 4032 7644
rect 3656 7590 3658 7642
rect 3658 7590 3710 7642
rect 3710 7590 3712 7642
rect 3736 7590 3774 7642
rect 3774 7590 3786 7642
rect 3786 7590 3792 7642
rect 3816 7590 3838 7642
rect 3838 7590 3850 7642
rect 3850 7590 3872 7642
rect 3896 7590 3902 7642
rect 3902 7590 3914 7642
rect 3914 7590 3952 7642
rect 3976 7590 3978 7642
rect 3978 7590 4030 7642
rect 4030 7590 4032 7642
rect 3656 7588 3712 7590
rect 3736 7588 3792 7590
rect 3816 7588 3872 7590
rect 3896 7588 3952 7590
rect 3976 7588 4032 7590
rect 2916 7098 2972 7100
rect 2996 7098 3052 7100
rect 3076 7098 3132 7100
rect 3156 7098 3212 7100
rect 3236 7098 3292 7100
rect 2916 7046 2918 7098
rect 2918 7046 2970 7098
rect 2970 7046 2972 7098
rect 2996 7046 3034 7098
rect 3034 7046 3046 7098
rect 3046 7046 3052 7098
rect 3076 7046 3098 7098
rect 3098 7046 3110 7098
rect 3110 7046 3132 7098
rect 3156 7046 3162 7098
rect 3162 7046 3174 7098
rect 3174 7046 3212 7098
rect 3236 7046 3238 7098
rect 3238 7046 3290 7098
rect 3290 7046 3292 7098
rect 2916 7044 2972 7046
rect 2996 7044 3052 7046
rect 3076 7044 3132 7046
rect 3156 7044 3212 7046
rect 3236 7044 3292 7046
rect 3606 7384 3662 7440
rect 3656 6554 3712 6556
rect 3736 6554 3792 6556
rect 3816 6554 3872 6556
rect 3896 6554 3952 6556
rect 3976 6554 4032 6556
rect 3656 6502 3658 6554
rect 3658 6502 3710 6554
rect 3710 6502 3712 6554
rect 3736 6502 3774 6554
rect 3774 6502 3786 6554
rect 3786 6502 3792 6554
rect 3816 6502 3838 6554
rect 3838 6502 3850 6554
rect 3850 6502 3872 6554
rect 3896 6502 3902 6554
rect 3902 6502 3914 6554
rect 3914 6502 3952 6554
rect 3976 6502 3978 6554
rect 3978 6502 4030 6554
rect 4030 6502 4032 6554
rect 3656 6500 3712 6502
rect 3736 6500 3792 6502
rect 3816 6500 3872 6502
rect 3896 6500 3952 6502
rect 3976 6500 4032 6502
rect 2916 6010 2972 6012
rect 2996 6010 3052 6012
rect 3076 6010 3132 6012
rect 3156 6010 3212 6012
rect 3236 6010 3292 6012
rect 2916 5958 2918 6010
rect 2918 5958 2970 6010
rect 2970 5958 2972 6010
rect 2996 5958 3034 6010
rect 3034 5958 3046 6010
rect 3046 5958 3052 6010
rect 3076 5958 3098 6010
rect 3098 5958 3110 6010
rect 3110 5958 3132 6010
rect 3156 5958 3162 6010
rect 3162 5958 3174 6010
rect 3174 5958 3212 6010
rect 3236 5958 3238 6010
rect 3238 5958 3290 6010
rect 3290 5958 3292 6010
rect 2916 5956 2972 5958
rect 2996 5956 3052 5958
rect 3076 5956 3132 5958
rect 3156 5956 3212 5958
rect 3236 5956 3292 5958
rect 3656 5466 3712 5468
rect 3736 5466 3792 5468
rect 3816 5466 3872 5468
rect 3896 5466 3952 5468
rect 3976 5466 4032 5468
rect 3656 5414 3658 5466
rect 3658 5414 3710 5466
rect 3710 5414 3712 5466
rect 3736 5414 3774 5466
rect 3774 5414 3786 5466
rect 3786 5414 3792 5466
rect 3816 5414 3838 5466
rect 3838 5414 3850 5466
rect 3850 5414 3872 5466
rect 3896 5414 3902 5466
rect 3902 5414 3914 5466
rect 3914 5414 3952 5466
rect 3976 5414 3978 5466
rect 3978 5414 4030 5466
rect 4030 5414 4032 5466
rect 3656 5412 3712 5414
rect 3736 5412 3792 5414
rect 3816 5412 3872 5414
rect 3896 5412 3952 5414
rect 3976 5412 4032 5414
rect 2916 4922 2972 4924
rect 2996 4922 3052 4924
rect 3076 4922 3132 4924
rect 3156 4922 3212 4924
rect 3236 4922 3292 4924
rect 2916 4870 2918 4922
rect 2918 4870 2970 4922
rect 2970 4870 2972 4922
rect 2996 4870 3034 4922
rect 3034 4870 3046 4922
rect 3046 4870 3052 4922
rect 3076 4870 3098 4922
rect 3098 4870 3110 4922
rect 3110 4870 3132 4922
rect 3156 4870 3162 4922
rect 3162 4870 3174 4922
rect 3174 4870 3212 4922
rect 3236 4870 3238 4922
rect 3238 4870 3290 4922
rect 3290 4870 3292 4922
rect 2916 4868 2972 4870
rect 2996 4868 3052 4870
rect 3076 4868 3132 4870
rect 3156 4868 3212 4870
rect 3236 4868 3292 4870
rect 3656 4378 3712 4380
rect 3736 4378 3792 4380
rect 3816 4378 3872 4380
rect 3896 4378 3952 4380
rect 3976 4378 4032 4380
rect 3656 4326 3658 4378
rect 3658 4326 3710 4378
rect 3710 4326 3712 4378
rect 3736 4326 3774 4378
rect 3774 4326 3786 4378
rect 3786 4326 3792 4378
rect 3816 4326 3838 4378
rect 3838 4326 3850 4378
rect 3850 4326 3872 4378
rect 3896 4326 3902 4378
rect 3902 4326 3914 4378
rect 3914 4326 3952 4378
rect 3976 4326 3978 4378
rect 3978 4326 4030 4378
rect 4030 4326 4032 4378
rect 3656 4324 3712 4326
rect 3736 4324 3792 4326
rect 3816 4324 3872 4326
rect 3896 4324 3952 4326
rect 3976 4324 4032 4326
rect 2916 3834 2972 3836
rect 2996 3834 3052 3836
rect 3076 3834 3132 3836
rect 3156 3834 3212 3836
rect 3236 3834 3292 3836
rect 2916 3782 2918 3834
rect 2918 3782 2970 3834
rect 2970 3782 2972 3834
rect 2996 3782 3034 3834
rect 3034 3782 3046 3834
rect 3046 3782 3052 3834
rect 3076 3782 3098 3834
rect 3098 3782 3110 3834
rect 3110 3782 3132 3834
rect 3156 3782 3162 3834
rect 3162 3782 3174 3834
rect 3174 3782 3212 3834
rect 3236 3782 3238 3834
rect 3238 3782 3290 3834
rect 3290 3782 3292 3834
rect 2916 3780 2972 3782
rect 2996 3780 3052 3782
rect 3076 3780 3132 3782
rect 3156 3780 3212 3782
rect 3236 3780 3292 3782
rect 3656 3290 3712 3292
rect 3736 3290 3792 3292
rect 3816 3290 3872 3292
rect 3896 3290 3952 3292
rect 3976 3290 4032 3292
rect 3656 3238 3658 3290
rect 3658 3238 3710 3290
rect 3710 3238 3712 3290
rect 3736 3238 3774 3290
rect 3774 3238 3786 3290
rect 3786 3238 3792 3290
rect 3816 3238 3838 3290
rect 3838 3238 3850 3290
rect 3850 3238 3872 3290
rect 3896 3238 3902 3290
rect 3902 3238 3914 3290
rect 3914 3238 3952 3290
rect 3976 3238 3978 3290
rect 3978 3238 4030 3290
rect 4030 3238 4032 3290
rect 3656 3236 3712 3238
rect 3736 3236 3792 3238
rect 3816 3236 3872 3238
rect 3896 3236 3952 3238
rect 3976 3236 4032 3238
rect 5170 8508 5172 8528
rect 5172 8508 5224 8528
rect 5224 8508 5226 8528
rect 5170 8472 5226 8508
rect 4526 7384 4582 7440
rect 5170 6996 5226 7032
rect 5170 6976 5172 6996
rect 5172 6976 5224 6996
rect 5224 6976 5226 6996
rect 5722 7384 5778 7440
rect 6916 21242 6972 21244
rect 6996 21242 7052 21244
rect 7076 21242 7132 21244
rect 7156 21242 7212 21244
rect 7236 21242 7292 21244
rect 6916 21190 6918 21242
rect 6918 21190 6970 21242
rect 6970 21190 6972 21242
rect 6996 21190 7034 21242
rect 7034 21190 7046 21242
rect 7046 21190 7052 21242
rect 7076 21190 7098 21242
rect 7098 21190 7110 21242
rect 7110 21190 7132 21242
rect 7156 21190 7162 21242
rect 7162 21190 7174 21242
rect 7174 21190 7212 21242
rect 7236 21190 7238 21242
rect 7238 21190 7290 21242
rect 7290 21190 7292 21242
rect 6916 21188 6972 21190
rect 6996 21188 7052 21190
rect 7076 21188 7132 21190
rect 7156 21188 7212 21190
rect 7236 21188 7292 21190
rect 6916 20154 6972 20156
rect 6996 20154 7052 20156
rect 7076 20154 7132 20156
rect 7156 20154 7212 20156
rect 7236 20154 7292 20156
rect 6916 20102 6918 20154
rect 6918 20102 6970 20154
rect 6970 20102 6972 20154
rect 6996 20102 7034 20154
rect 7034 20102 7046 20154
rect 7046 20102 7052 20154
rect 7076 20102 7098 20154
rect 7098 20102 7110 20154
rect 7110 20102 7132 20154
rect 7156 20102 7162 20154
rect 7162 20102 7174 20154
rect 7174 20102 7212 20154
rect 7236 20102 7238 20154
rect 7238 20102 7290 20154
rect 7290 20102 7292 20154
rect 6916 20100 6972 20102
rect 6996 20100 7052 20102
rect 7076 20100 7132 20102
rect 7156 20100 7212 20102
rect 7236 20100 7292 20102
rect 7656 22874 7712 22876
rect 7736 22874 7792 22876
rect 7816 22874 7872 22876
rect 7896 22874 7952 22876
rect 7976 22874 8032 22876
rect 7656 22822 7658 22874
rect 7658 22822 7710 22874
rect 7710 22822 7712 22874
rect 7736 22822 7774 22874
rect 7774 22822 7786 22874
rect 7786 22822 7792 22874
rect 7816 22822 7838 22874
rect 7838 22822 7850 22874
rect 7850 22822 7872 22874
rect 7896 22822 7902 22874
rect 7902 22822 7914 22874
rect 7914 22822 7952 22874
rect 7976 22822 7978 22874
rect 7978 22822 8030 22874
rect 8030 22822 8032 22874
rect 7656 22820 7712 22822
rect 7736 22820 7792 22822
rect 7816 22820 7872 22822
rect 7896 22820 7952 22822
rect 7976 22820 8032 22822
rect 7656 21786 7712 21788
rect 7736 21786 7792 21788
rect 7816 21786 7872 21788
rect 7896 21786 7952 21788
rect 7976 21786 8032 21788
rect 7656 21734 7658 21786
rect 7658 21734 7710 21786
rect 7710 21734 7712 21786
rect 7736 21734 7774 21786
rect 7774 21734 7786 21786
rect 7786 21734 7792 21786
rect 7816 21734 7838 21786
rect 7838 21734 7850 21786
rect 7850 21734 7872 21786
rect 7896 21734 7902 21786
rect 7902 21734 7914 21786
rect 7914 21734 7952 21786
rect 7976 21734 7978 21786
rect 7978 21734 8030 21786
rect 8030 21734 8032 21786
rect 7656 21732 7712 21734
rect 7736 21732 7792 21734
rect 7816 21732 7872 21734
rect 7896 21732 7952 21734
rect 7976 21732 8032 21734
rect 7656 20698 7712 20700
rect 7736 20698 7792 20700
rect 7816 20698 7872 20700
rect 7896 20698 7952 20700
rect 7976 20698 8032 20700
rect 7656 20646 7658 20698
rect 7658 20646 7710 20698
rect 7710 20646 7712 20698
rect 7736 20646 7774 20698
rect 7774 20646 7786 20698
rect 7786 20646 7792 20698
rect 7816 20646 7838 20698
rect 7838 20646 7850 20698
rect 7850 20646 7872 20698
rect 7896 20646 7902 20698
rect 7902 20646 7914 20698
rect 7914 20646 7952 20698
rect 7976 20646 7978 20698
rect 7978 20646 8030 20698
rect 8030 20646 8032 20698
rect 7656 20644 7712 20646
rect 7736 20644 7792 20646
rect 7816 20644 7872 20646
rect 7896 20644 7952 20646
rect 7976 20644 8032 20646
rect 7656 19610 7712 19612
rect 7736 19610 7792 19612
rect 7816 19610 7872 19612
rect 7896 19610 7952 19612
rect 7976 19610 8032 19612
rect 7656 19558 7658 19610
rect 7658 19558 7710 19610
rect 7710 19558 7712 19610
rect 7736 19558 7774 19610
rect 7774 19558 7786 19610
rect 7786 19558 7792 19610
rect 7816 19558 7838 19610
rect 7838 19558 7850 19610
rect 7850 19558 7872 19610
rect 7896 19558 7902 19610
rect 7902 19558 7914 19610
rect 7914 19558 7952 19610
rect 7976 19558 7978 19610
rect 7978 19558 8030 19610
rect 8030 19558 8032 19610
rect 7656 19556 7712 19558
rect 7736 19556 7792 19558
rect 7816 19556 7872 19558
rect 7896 19556 7952 19558
rect 7976 19556 8032 19558
rect 6916 19066 6972 19068
rect 6996 19066 7052 19068
rect 7076 19066 7132 19068
rect 7156 19066 7212 19068
rect 7236 19066 7292 19068
rect 6916 19014 6918 19066
rect 6918 19014 6970 19066
rect 6970 19014 6972 19066
rect 6996 19014 7034 19066
rect 7034 19014 7046 19066
rect 7046 19014 7052 19066
rect 7076 19014 7098 19066
rect 7098 19014 7110 19066
rect 7110 19014 7132 19066
rect 7156 19014 7162 19066
rect 7162 19014 7174 19066
rect 7174 19014 7212 19066
rect 7236 19014 7238 19066
rect 7238 19014 7290 19066
rect 7290 19014 7292 19066
rect 6916 19012 6972 19014
rect 6996 19012 7052 19014
rect 7076 19012 7132 19014
rect 7156 19012 7212 19014
rect 7236 19012 7292 19014
rect 6916 17978 6972 17980
rect 6996 17978 7052 17980
rect 7076 17978 7132 17980
rect 7156 17978 7212 17980
rect 7236 17978 7292 17980
rect 6916 17926 6918 17978
rect 6918 17926 6970 17978
rect 6970 17926 6972 17978
rect 6996 17926 7034 17978
rect 7034 17926 7046 17978
rect 7046 17926 7052 17978
rect 7076 17926 7098 17978
rect 7098 17926 7110 17978
rect 7110 17926 7132 17978
rect 7156 17926 7162 17978
rect 7162 17926 7174 17978
rect 7174 17926 7212 17978
rect 7236 17926 7238 17978
rect 7238 17926 7290 17978
rect 7290 17926 7292 17978
rect 6916 17924 6972 17926
rect 6996 17924 7052 17926
rect 7076 17924 7132 17926
rect 7156 17924 7212 17926
rect 7236 17924 7292 17926
rect 6916 16890 6972 16892
rect 6996 16890 7052 16892
rect 7076 16890 7132 16892
rect 7156 16890 7212 16892
rect 7236 16890 7292 16892
rect 6916 16838 6918 16890
rect 6918 16838 6970 16890
rect 6970 16838 6972 16890
rect 6996 16838 7034 16890
rect 7034 16838 7046 16890
rect 7046 16838 7052 16890
rect 7076 16838 7098 16890
rect 7098 16838 7110 16890
rect 7110 16838 7132 16890
rect 7156 16838 7162 16890
rect 7162 16838 7174 16890
rect 7174 16838 7212 16890
rect 7236 16838 7238 16890
rect 7238 16838 7290 16890
rect 7290 16838 7292 16890
rect 6916 16836 6972 16838
rect 6996 16836 7052 16838
rect 7076 16836 7132 16838
rect 7156 16836 7212 16838
rect 7236 16836 7292 16838
rect 6916 15802 6972 15804
rect 6996 15802 7052 15804
rect 7076 15802 7132 15804
rect 7156 15802 7212 15804
rect 7236 15802 7292 15804
rect 6916 15750 6918 15802
rect 6918 15750 6970 15802
rect 6970 15750 6972 15802
rect 6996 15750 7034 15802
rect 7034 15750 7046 15802
rect 7046 15750 7052 15802
rect 7076 15750 7098 15802
rect 7098 15750 7110 15802
rect 7110 15750 7132 15802
rect 7156 15750 7162 15802
rect 7162 15750 7174 15802
rect 7174 15750 7212 15802
rect 7236 15750 7238 15802
rect 7238 15750 7290 15802
rect 7290 15750 7292 15802
rect 6916 15748 6972 15750
rect 6996 15748 7052 15750
rect 7076 15748 7132 15750
rect 7156 15748 7212 15750
rect 7236 15748 7292 15750
rect 7656 18522 7712 18524
rect 7736 18522 7792 18524
rect 7816 18522 7872 18524
rect 7896 18522 7952 18524
rect 7976 18522 8032 18524
rect 7656 18470 7658 18522
rect 7658 18470 7710 18522
rect 7710 18470 7712 18522
rect 7736 18470 7774 18522
rect 7774 18470 7786 18522
rect 7786 18470 7792 18522
rect 7816 18470 7838 18522
rect 7838 18470 7850 18522
rect 7850 18470 7872 18522
rect 7896 18470 7902 18522
rect 7902 18470 7914 18522
rect 7914 18470 7952 18522
rect 7976 18470 7978 18522
rect 7978 18470 8030 18522
rect 8030 18470 8032 18522
rect 7656 18468 7712 18470
rect 7736 18468 7792 18470
rect 7816 18468 7872 18470
rect 7896 18468 7952 18470
rect 7976 18468 8032 18470
rect 7656 17434 7712 17436
rect 7736 17434 7792 17436
rect 7816 17434 7872 17436
rect 7896 17434 7952 17436
rect 7976 17434 8032 17436
rect 7656 17382 7658 17434
rect 7658 17382 7710 17434
rect 7710 17382 7712 17434
rect 7736 17382 7774 17434
rect 7774 17382 7786 17434
rect 7786 17382 7792 17434
rect 7816 17382 7838 17434
rect 7838 17382 7850 17434
rect 7850 17382 7872 17434
rect 7896 17382 7902 17434
rect 7902 17382 7914 17434
rect 7914 17382 7952 17434
rect 7976 17382 7978 17434
rect 7978 17382 8030 17434
rect 8030 17382 8032 17434
rect 7656 17380 7712 17382
rect 7736 17380 7792 17382
rect 7816 17380 7872 17382
rect 7896 17380 7952 17382
rect 7976 17380 8032 17382
rect 7656 16346 7712 16348
rect 7736 16346 7792 16348
rect 7816 16346 7872 16348
rect 7896 16346 7952 16348
rect 7976 16346 8032 16348
rect 7656 16294 7658 16346
rect 7658 16294 7710 16346
rect 7710 16294 7712 16346
rect 7736 16294 7774 16346
rect 7774 16294 7786 16346
rect 7786 16294 7792 16346
rect 7816 16294 7838 16346
rect 7838 16294 7850 16346
rect 7850 16294 7872 16346
rect 7896 16294 7902 16346
rect 7902 16294 7914 16346
rect 7914 16294 7952 16346
rect 7976 16294 7978 16346
rect 7978 16294 8030 16346
rect 8030 16294 8032 16346
rect 7656 16292 7712 16294
rect 7736 16292 7792 16294
rect 7816 16292 7872 16294
rect 7896 16292 7952 16294
rect 7976 16292 8032 16294
rect 6916 14714 6972 14716
rect 6996 14714 7052 14716
rect 7076 14714 7132 14716
rect 7156 14714 7212 14716
rect 7236 14714 7292 14716
rect 6916 14662 6918 14714
rect 6918 14662 6970 14714
rect 6970 14662 6972 14714
rect 6996 14662 7034 14714
rect 7034 14662 7046 14714
rect 7046 14662 7052 14714
rect 7076 14662 7098 14714
rect 7098 14662 7110 14714
rect 7110 14662 7132 14714
rect 7156 14662 7162 14714
rect 7162 14662 7174 14714
rect 7174 14662 7212 14714
rect 7236 14662 7238 14714
rect 7238 14662 7290 14714
rect 7290 14662 7292 14714
rect 6916 14660 6972 14662
rect 6996 14660 7052 14662
rect 7076 14660 7132 14662
rect 7156 14660 7212 14662
rect 7236 14660 7292 14662
rect 7656 15258 7712 15260
rect 7736 15258 7792 15260
rect 7816 15258 7872 15260
rect 7896 15258 7952 15260
rect 7976 15258 8032 15260
rect 7656 15206 7658 15258
rect 7658 15206 7710 15258
rect 7710 15206 7712 15258
rect 7736 15206 7774 15258
rect 7774 15206 7786 15258
rect 7786 15206 7792 15258
rect 7816 15206 7838 15258
rect 7838 15206 7850 15258
rect 7850 15206 7872 15258
rect 7896 15206 7902 15258
rect 7902 15206 7914 15258
rect 7914 15206 7952 15258
rect 7976 15206 7978 15258
rect 7978 15206 8030 15258
rect 8030 15206 8032 15258
rect 7656 15204 7712 15206
rect 7736 15204 7792 15206
rect 7816 15204 7872 15206
rect 7896 15204 7952 15206
rect 7976 15204 8032 15206
rect 7746 14864 7802 14920
rect 7656 14170 7712 14172
rect 7736 14170 7792 14172
rect 7816 14170 7872 14172
rect 7896 14170 7952 14172
rect 7976 14170 8032 14172
rect 7656 14118 7658 14170
rect 7658 14118 7710 14170
rect 7710 14118 7712 14170
rect 7736 14118 7774 14170
rect 7774 14118 7786 14170
rect 7786 14118 7792 14170
rect 7816 14118 7838 14170
rect 7838 14118 7850 14170
rect 7850 14118 7872 14170
rect 7896 14118 7902 14170
rect 7902 14118 7914 14170
rect 7914 14118 7952 14170
rect 7976 14118 7978 14170
rect 7978 14118 8030 14170
rect 8030 14118 8032 14170
rect 7656 14116 7712 14118
rect 7736 14116 7792 14118
rect 7816 14116 7872 14118
rect 7896 14116 7952 14118
rect 7976 14116 8032 14118
rect 6916 13626 6972 13628
rect 6996 13626 7052 13628
rect 7076 13626 7132 13628
rect 7156 13626 7212 13628
rect 7236 13626 7292 13628
rect 6916 13574 6918 13626
rect 6918 13574 6970 13626
rect 6970 13574 6972 13626
rect 6996 13574 7034 13626
rect 7034 13574 7046 13626
rect 7046 13574 7052 13626
rect 7076 13574 7098 13626
rect 7098 13574 7110 13626
rect 7110 13574 7132 13626
rect 7156 13574 7162 13626
rect 7162 13574 7174 13626
rect 7174 13574 7212 13626
rect 7236 13574 7238 13626
rect 7238 13574 7290 13626
rect 7290 13574 7292 13626
rect 6916 13572 6972 13574
rect 6996 13572 7052 13574
rect 7076 13572 7132 13574
rect 7156 13572 7212 13574
rect 7236 13572 7292 13574
rect 6916 12538 6972 12540
rect 6996 12538 7052 12540
rect 7076 12538 7132 12540
rect 7156 12538 7212 12540
rect 7236 12538 7292 12540
rect 6916 12486 6918 12538
rect 6918 12486 6970 12538
rect 6970 12486 6972 12538
rect 6996 12486 7034 12538
rect 7034 12486 7046 12538
rect 7046 12486 7052 12538
rect 7076 12486 7098 12538
rect 7098 12486 7110 12538
rect 7110 12486 7132 12538
rect 7156 12486 7162 12538
rect 7162 12486 7174 12538
rect 7174 12486 7212 12538
rect 7236 12486 7238 12538
rect 7238 12486 7290 12538
rect 7290 12486 7292 12538
rect 6916 12484 6972 12486
rect 6996 12484 7052 12486
rect 7076 12484 7132 12486
rect 7156 12484 7212 12486
rect 7236 12484 7292 12486
rect 7656 13082 7712 13084
rect 7736 13082 7792 13084
rect 7816 13082 7872 13084
rect 7896 13082 7952 13084
rect 7976 13082 8032 13084
rect 7656 13030 7658 13082
rect 7658 13030 7710 13082
rect 7710 13030 7712 13082
rect 7736 13030 7774 13082
rect 7774 13030 7786 13082
rect 7786 13030 7792 13082
rect 7816 13030 7838 13082
rect 7838 13030 7850 13082
rect 7850 13030 7872 13082
rect 7896 13030 7902 13082
rect 7902 13030 7914 13082
rect 7914 13030 7952 13082
rect 7976 13030 7978 13082
rect 7978 13030 8030 13082
rect 8030 13030 8032 13082
rect 7656 13028 7712 13030
rect 7736 13028 7792 13030
rect 7816 13028 7872 13030
rect 7896 13028 7952 13030
rect 7976 13028 8032 13030
rect 6916 11450 6972 11452
rect 6996 11450 7052 11452
rect 7076 11450 7132 11452
rect 7156 11450 7212 11452
rect 7236 11450 7292 11452
rect 6916 11398 6918 11450
rect 6918 11398 6970 11450
rect 6970 11398 6972 11450
rect 6996 11398 7034 11450
rect 7034 11398 7046 11450
rect 7046 11398 7052 11450
rect 7076 11398 7098 11450
rect 7098 11398 7110 11450
rect 7110 11398 7132 11450
rect 7156 11398 7162 11450
rect 7162 11398 7174 11450
rect 7174 11398 7212 11450
rect 7236 11398 7238 11450
rect 7238 11398 7290 11450
rect 7290 11398 7292 11450
rect 6916 11396 6972 11398
rect 6996 11396 7052 11398
rect 7076 11396 7132 11398
rect 7156 11396 7212 11398
rect 7236 11396 7292 11398
rect 7656 11994 7712 11996
rect 7736 11994 7792 11996
rect 7816 11994 7872 11996
rect 7896 11994 7952 11996
rect 7976 11994 8032 11996
rect 7656 11942 7658 11994
rect 7658 11942 7710 11994
rect 7710 11942 7712 11994
rect 7736 11942 7774 11994
rect 7774 11942 7786 11994
rect 7786 11942 7792 11994
rect 7816 11942 7838 11994
rect 7838 11942 7850 11994
rect 7850 11942 7872 11994
rect 7896 11942 7902 11994
rect 7902 11942 7914 11994
rect 7914 11942 7952 11994
rect 7976 11942 7978 11994
rect 7978 11942 8030 11994
rect 8030 11942 8032 11994
rect 7656 11940 7712 11942
rect 7736 11940 7792 11942
rect 7816 11940 7872 11942
rect 7896 11940 7952 11942
rect 7976 11940 8032 11942
rect 7656 10906 7712 10908
rect 7736 10906 7792 10908
rect 7816 10906 7872 10908
rect 7896 10906 7952 10908
rect 7976 10906 8032 10908
rect 7656 10854 7658 10906
rect 7658 10854 7710 10906
rect 7710 10854 7712 10906
rect 7736 10854 7774 10906
rect 7774 10854 7786 10906
rect 7786 10854 7792 10906
rect 7816 10854 7838 10906
rect 7838 10854 7850 10906
rect 7850 10854 7872 10906
rect 7896 10854 7902 10906
rect 7902 10854 7914 10906
rect 7914 10854 7952 10906
rect 7976 10854 7978 10906
rect 7978 10854 8030 10906
rect 8030 10854 8032 10906
rect 7656 10852 7712 10854
rect 7736 10852 7792 10854
rect 7816 10852 7872 10854
rect 7896 10852 7952 10854
rect 7976 10852 8032 10854
rect 6916 10362 6972 10364
rect 6996 10362 7052 10364
rect 7076 10362 7132 10364
rect 7156 10362 7212 10364
rect 7236 10362 7292 10364
rect 6916 10310 6918 10362
rect 6918 10310 6970 10362
rect 6970 10310 6972 10362
rect 6996 10310 7034 10362
rect 7034 10310 7046 10362
rect 7046 10310 7052 10362
rect 7076 10310 7098 10362
rect 7098 10310 7110 10362
rect 7110 10310 7132 10362
rect 7156 10310 7162 10362
rect 7162 10310 7174 10362
rect 7174 10310 7212 10362
rect 7236 10310 7238 10362
rect 7238 10310 7290 10362
rect 7290 10310 7292 10362
rect 6916 10308 6972 10310
rect 6996 10308 7052 10310
rect 7076 10308 7132 10310
rect 7156 10308 7212 10310
rect 7236 10308 7292 10310
rect 7102 10124 7158 10160
rect 7102 10104 7104 10124
rect 7104 10104 7156 10124
rect 7156 10104 7158 10124
rect 8114 10512 8170 10568
rect 7562 10260 7618 10296
rect 7562 10240 7564 10260
rect 7564 10240 7616 10260
rect 7616 10240 7618 10260
rect 8298 10512 8354 10568
rect 7656 9818 7712 9820
rect 7736 9818 7792 9820
rect 7816 9818 7872 9820
rect 7896 9818 7952 9820
rect 7976 9818 8032 9820
rect 7656 9766 7658 9818
rect 7658 9766 7710 9818
rect 7710 9766 7712 9818
rect 7736 9766 7774 9818
rect 7774 9766 7786 9818
rect 7786 9766 7792 9818
rect 7816 9766 7838 9818
rect 7838 9766 7850 9818
rect 7850 9766 7872 9818
rect 7896 9766 7902 9818
rect 7902 9766 7914 9818
rect 7914 9766 7952 9818
rect 7976 9766 7978 9818
rect 7978 9766 8030 9818
rect 8030 9766 8032 9818
rect 7656 9764 7712 9766
rect 7736 9764 7792 9766
rect 7816 9764 7872 9766
rect 7896 9764 7952 9766
rect 7976 9764 8032 9766
rect 6916 9274 6972 9276
rect 6996 9274 7052 9276
rect 7076 9274 7132 9276
rect 7156 9274 7212 9276
rect 7236 9274 7292 9276
rect 6916 9222 6918 9274
rect 6918 9222 6970 9274
rect 6970 9222 6972 9274
rect 6996 9222 7034 9274
rect 7034 9222 7046 9274
rect 7046 9222 7052 9274
rect 7076 9222 7098 9274
rect 7098 9222 7110 9274
rect 7110 9222 7132 9274
rect 7156 9222 7162 9274
rect 7162 9222 7174 9274
rect 7174 9222 7212 9274
rect 7236 9222 7238 9274
rect 7238 9222 7290 9274
rect 7290 9222 7292 9274
rect 6916 9220 6972 9222
rect 6996 9220 7052 9222
rect 7076 9220 7132 9222
rect 7156 9220 7212 9222
rect 7236 9220 7292 9222
rect 7656 8730 7712 8732
rect 7736 8730 7792 8732
rect 7816 8730 7872 8732
rect 7896 8730 7952 8732
rect 7976 8730 8032 8732
rect 7656 8678 7658 8730
rect 7658 8678 7710 8730
rect 7710 8678 7712 8730
rect 7736 8678 7774 8730
rect 7774 8678 7786 8730
rect 7786 8678 7792 8730
rect 7816 8678 7838 8730
rect 7838 8678 7850 8730
rect 7850 8678 7872 8730
rect 7896 8678 7902 8730
rect 7902 8678 7914 8730
rect 7914 8678 7952 8730
rect 7976 8678 7978 8730
rect 7978 8678 8030 8730
rect 8030 8678 8032 8730
rect 7656 8676 7712 8678
rect 7736 8676 7792 8678
rect 7816 8676 7872 8678
rect 7896 8676 7952 8678
rect 7976 8676 8032 8678
rect 6916 8186 6972 8188
rect 6996 8186 7052 8188
rect 7076 8186 7132 8188
rect 7156 8186 7212 8188
rect 7236 8186 7292 8188
rect 6916 8134 6918 8186
rect 6918 8134 6970 8186
rect 6970 8134 6972 8186
rect 6996 8134 7034 8186
rect 7034 8134 7046 8186
rect 7046 8134 7052 8186
rect 7076 8134 7098 8186
rect 7098 8134 7110 8186
rect 7110 8134 7132 8186
rect 7156 8134 7162 8186
rect 7162 8134 7174 8186
rect 7174 8134 7212 8186
rect 7236 8134 7238 8186
rect 7238 8134 7290 8186
rect 7290 8134 7292 8186
rect 6916 8132 6972 8134
rect 6996 8132 7052 8134
rect 7076 8132 7132 8134
rect 7156 8132 7212 8134
rect 7236 8132 7292 8134
rect 8482 9968 8538 10024
rect 7656 7642 7712 7644
rect 7736 7642 7792 7644
rect 7816 7642 7872 7644
rect 7896 7642 7952 7644
rect 7976 7642 8032 7644
rect 7656 7590 7658 7642
rect 7658 7590 7710 7642
rect 7710 7590 7712 7642
rect 7736 7590 7774 7642
rect 7774 7590 7786 7642
rect 7786 7590 7792 7642
rect 7816 7590 7838 7642
rect 7838 7590 7850 7642
rect 7850 7590 7872 7642
rect 7896 7590 7902 7642
rect 7902 7590 7914 7642
rect 7914 7590 7952 7642
rect 7976 7590 7978 7642
rect 7978 7590 8030 7642
rect 8030 7590 8032 7642
rect 7656 7588 7712 7590
rect 7736 7588 7792 7590
rect 7816 7588 7872 7590
rect 7896 7588 7952 7590
rect 7976 7588 8032 7590
rect 6916 7098 6972 7100
rect 6996 7098 7052 7100
rect 7076 7098 7132 7100
rect 7156 7098 7212 7100
rect 7236 7098 7292 7100
rect 6916 7046 6918 7098
rect 6918 7046 6970 7098
rect 6970 7046 6972 7098
rect 6996 7046 7034 7098
rect 7034 7046 7046 7098
rect 7046 7046 7052 7098
rect 7076 7046 7098 7098
rect 7098 7046 7110 7098
rect 7110 7046 7132 7098
rect 7156 7046 7162 7098
rect 7162 7046 7174 7098
rect 7174 7046 7212 7098
rect 7236 7046 7238 7098
rect 7238 7046 7290 7098
rect 7290 7046 7292 7098
rect 6916 7044 6972 7046
rect 6996 7044 7052 7046
rect 7076 7044 7132 7046
rect 7156 7044 7212 7046
rect 7236 7044 7292 7046
rect 6916 6010 6972 6012
rect 6996 6010 7052 6012
rect 7076 6010 7132 6012
rect 7156 6010 7212 6012
rect 7236 6010 7292 6012
rect 6916 5958 6918 6010
rect 6918 5958 6970 6010
rect 6970 5958 6972 6010
rect 6996 5958 7034 6010
rect 7034 5958 7046 6010
rect 7046 5958 7052 6010
rect 7076 5958 7098 6010
rect 7098 5958 7110 6010
rect 7110 5958 7132 6010
rect 7156 5958 7162 6010
rect 7162 5958 7174 6010
rect 7174 5958 7212 6010
rect 7236 5958 7238 6010
rect 7238 5958 7290 6010
rect 7290 5958 7292 6010
rect 6916 5956 6972 5958
rect 6996 5956 7052 5958
rect 7076 5956 7132 5958
rect 7156 5956 7212 5958
rect 7236 5956 7292 5958
rect 7746 7384 7802 7440
rect 8298 7384 8354 7440
rect 7656 6554 7712 6556
rect 7736 6554 7792 6556
rect 7816 6554 7872 6556
rect 7896 6554 7952 6556
rect 7976 6554 8032 6556
rect 7656 6502 7658 6554
rect 7658 6502 7710 6554
rect 7710 6502 7712 6554
rect 7736 6502 7774 6554
rect 7774 6502 7786 6554
rect 7786 6502 7792 6554
rect 7816 6502 7838 6554
rect 7838 6502 7850 6554
rect 7850 6502 7872 6554
rect 7896 6502 7902 6554
rect 7902 6502 7914 6554
rect 7914 6502 7952 6554
rect 7976 6502 7978 6554
rect 7978 6502 8030 6554
rect 8030 6502 8032 6554
rect 7656 6500 7712 6502
rect 7736 6500 7792 6502
rect 7816 6500 7872 6502
rect 7896 6500 7952 6502
rect 7976 6500 8032 6502
rect 6916 4922 6972 4924
rect 6996 4922 7052 4924
rect 7076 4922 7132 4924
rect 7156 4922 7212 4924
rect 7236 4922 7292 4924
rect 6916 4870 6918 4922
rect 6918 4870 6970 4922
rect 6970 4870 6972 4922
rect 6996 4870 7034 4922
rect 7034 4870 7046 4922
rect 7046 4870 7052 4922
rect 7076 4870 7098 4922
rect 7098 4870 7110 4922
rect 7110 4870 7132 4922
rect 7156 4870 7162 4922
rect 7162 4870 7174 4922
rect 7174 4870 7212 4922
rect 7236 4870 7238 4922
rect 7238 4870 7290 4922
rect 7290 4870 7292 4922
rect 6916 4868 6972 4870
rect 6996 4868 7052 4870
rect 7076 4868 7132 4870
rect 7156 4868 7212 4870
rect 7236 4868 7292 4870
rect 6916 3834 6972 3836
rect 6996 3834 7052 3836
rect 7076 3834 7132 3836
rect 7156 3834 7212 3836
rect 7236 3834 7292 3836
rect 6916 3782 6918 3834
rect 6918 3782 6970 3834
rect 6970 3782 6972 3834
rect 6996 3782 7034 3834
rect 7034 3782 7046 3834
rect 7046 3782 7052 3834
rect 7076 3782 7098 3834
rect 7098 3782 7110 3834
rect 7110 3782 7132 3834
rect 7156 3782 7162 3834
rect 7162 3782 7174 3834
rect 7174 3782 7212 3834
rect 7236 3782 7238 3834
rect 7238 3782 7290 3834
rect 7290 3782 7292 3834
rect 6916 3780 6972 3782
rect 6996 3780 7052 3782
rect 7076 3780 7132 3782
rect 7156 3780 7212 3782
rect 7236 3780 7292 3782
rect 2916 2746 2972 2748
rect 2996 2746 3052 2748
rect 3076 2746 3132 2748
rect 3156 2746 3212 2748
rect 3236 2746 3292 2748
rect 2916 2694 2918 2746
rect 2918 2694 2970 2746
rect 2970 2694 2972 2746
rect 2996 2694 3034 2746
rect 3034 2694 3046 2746
rect 3046 2694 3052 2746
rect 3076 2694 3098 2746
rect 3098 2694 3110 2746
rect 3110 2694 3132 2746
rect 3156 2694 3162 2746
rect 3162 2694 3174 2746
rect 3174 2694 3212 2746
rect 3236 2694 3238 2746
rect 3238 2694 3290 2746
rect 3290 2694 3292 2746
rect 2916 2692 2972 2694
rect 2996 2692 3052 2694
rect 3076 2692 3132 2694
rect 3156 2692 3212 2694
rect 3236 2692 3292 2694
rect 9126 15136 9182 15192
rect 9034 14864 9090 14920
rect 9678 18808 9734 18864
rect 9126 11736 9182 11792
rect 9034 10104 9090 10160
rect 9494 10240 9550 10296
rect 9586 9968 9642 10024
rect 10046 10804 10102 10840
rect 10874 26832 10930 26888
rect 10916 26682 10972 26684
rect 10996 26682 11052 26684
rect 11076 26682 11132 26684
rect 11156 26682 11212 26684
rect 11236 26682 11292 26684
rect 10916 26630 10918 26682
rect 10918 26630 10970 26682
rect 10970 26630 10972 26682
rect 10996 26630 11034 26682
rect 11034 26630 11046 26682
rect 11046 26630 11052 26682
rect 11076 26630 11098 26682
rect 11098 26630 11110 26682
rect 11110 26630 11132 26682
rect 11156 26630 11162 26682
rect 11162 26630 11174 26682
rect 11174 26630 11212 26682
rect 11236 26630 11238 26682
rect 11238 26630 11290 26682
rect 11290 26630 11292 26682
rect 10916 26628 10972 26630
rect 10996 26628 11052 26630
rect 11076 26628 11132 26630
rect 11156 26628 11212 26630
rect 11236 26628 11292 26630
rect 10916 25594 10972 25596
rect 10996 25594 11052 25596
rect 11076 25594 11132 25596
rect 11156 25594 11212 25596
rect 11236 25594 11292 25596
rect 10916 25542 10918 25594
rect 10918 25542 10970 25594
rect 10970 25542 10972 25594
rect 10996 25542 11034 25594
rect 11034 25542 11046 25594
rect 11046 25542 11052 25594
rect 11076 25542 11098 25594
rect 11098 25542 11110 25594
rect 11110 25542 11132 25594
rect 11156 25542 11162 25594
rect 11162 25542 11174 25594
rect 11174 25542 11212 25594
rect 11236 25542 11238 25594
rect 11238 25542 11290 25594
rect 11290 25542 11292 25594
rect 10916 25540 10972 25542
rect 10996 25540 11052 25542
rect 11076 25540 11132 25542
rect 11156 25540 11212 25542
rect 11236 25540 11292 25542
rect 10414 19372 10470 19408
rect 10414 19352 10416 19372
rect 10416 19352 10468 19372
rect 10468 19352 10470 19372
rect 10230 19252 10232 19272
rect 10232 19252 10284 19272
rect 10284 19252 10286 19272
rect 10230 19216 10286 19252
rect 10322 18808 10378 18864
rect 10414 18128 10470 18184
rect 10916 24506 10972 24508
rect 10996 24506 11052 24508
rect 11076 24506 11132 24508
rect 11156 24506 11212 24508
rect 11236 24506 11292 24508
rect 10916 24454 10918 24506
rect 10918 24454 10970 24506
rect 10970 24454 10972 24506
rect 10996 24454 11034 24506
rect 11034 24454 11046 24506
rect 11046 24454 11052 24506
rect 11076 24454 11098 24506
rect 11098 24454 11110 24506
rect 11110 24454 11132 24506
rect 11156 24454 11162 24506
rect 11162 24454 11174 24506
rect 11174 24454 11212 24506
rect 11236 24454 11238 24506
rect 11238 24454 11290 24506
rect 11290 24454 11292 24506
rect 10916 24452 10972 24454
rect 10996 24452 11052 24454
rect 11076 24452 11132 24454
rect 11156 24452 11212 24454
rect 11236 24452 11292 24454
rect 10916 23418 10972 23420
rect 10996 23418 11052 23420
rect 11076 23418 11132 23420
rect 11156 23418 11212 23420
rect 11236 23418 11292 23420
rect 10916 23366 10918 23418
rect 10918 23366 10970 23418
rect 10970 23366 10972 23418
rect 10996 23366 11034 23418
rect 11034 23366 11046 23418
rect 11046 23366 11052 23418
rect 11076 23366 11098 23418
rect 11098 23366 11110 23418
rect 11110 23366 11132 23418
rect 11156 23366 11162 23418
rect 11162 23366 11174 23418
rect 11174 23366 11212 23418
rect 11236 23366 11238 23418
rect 11238 23366 11290 23418
rect 11290 23366 11292 23418
rect 10916 23364 10972 23366
rect 10996 23364 11052 23366
rect 11076 23364 11132 23366
rect 11156 23364 11212 23366
rect 11236 23364 11292 23366
rect 10874 23024 10930 23080
rect 11656 27226 11712 27228
rect 11736 27226 11792 27228
rect 11816 27226 11872 27228
rect 11896 27226 11952 27228
rect 11976 27226 12032 27228
rect 11656 27174 11658 27226
rect 11658 27174 11710 27226
rect 11710 27174 11712 27226
rect 11736 27174 11774 27226
rect 11774 27174 11786 27226
rect 11786 27174 11792 27226
rect 11816 27174 11838 27226
rect 11838 27174 11850 27226
rect 11850 27174 11872 27226
rect 11896 27174 11902 27226
rect 11902 27174 11914 27226
rect 11914 27174 11952 27226
rect 11976 27174 11978 27226
rect 11978 27174 12030 27226
rect 12030 27174 12032 27226
rect 11656 27172 11712 27174
rect 11736 27172 11792 27174
rect 11816 27172 11872 27174
rect 11896 27172 11952 27174
rect 11976 27172 12032 27174
rect 11656 26138 11712 26140
rect 11736 26138 11792 26140
rect 11816 26138 11872 26140
rect 11896 26138 11952 26140
rect 11976 26138 12032 26140
rect 11656 26086 11658 26138
rect 11658 26086 11710 26138
rect 11710 26086 11712 26138
rect 11736 26086 11774 26138
rect 11774 26086 11786 26138
rect 11786 26086 11792 26138
rect 11816 26086 11838 26138
rect 11838 26086 11850 26138
rect 11850 26086 11872 26138
rect 11896 26086 11902 26138
rect 11902 26086 11914 26138
rect 11914 26086 11952 26138
rect 11976 26086 11978 26138
rect 11978 26086 12030 26138
rect 12030 26086 12032 26138
rect 11656 26084 11712 26086
rect 11736 26084 11792 26086
rect 11816 26084 11872 26086
rect 11896 26084 11952 26086
rect 11976 26084 12032 26086
rect 11656 25050 11712 25052
rect 11736 25050 11792 25052
rect 11816 25050 11872 25052
rect 11896 25050 11952 25052
rect 11976 25050 12032 25052
rect 11656 24998 11658 25050
rect 11658 24998 11710 25050
rect 11710 24998 11712 25050
rect 11736 24998 11774 25050
rect 11774 24998 11786 25050
rect 11786 24998 11792 25050
rect 11816 24998 11838 25050
rect 11838 24998 11850 25050
rect 11850 24998 11872 25050
rect 11896 24998 11902 25050
rect 11902 24998 11914 25050
rect 11914 24998 11952 25050
rect 11976 24998 11978 25050
rect 11978 24998 12030 25050
rect 12030 24998 12032 25050
rect 11656 24996 11712 24998
rect 11736 24996 11792 24998
rect 11816 24996 11872 24998
rect 11896 24996 11952 24998
rect 11976 24996 12032 24998
rect 11656 23962 11712 23964
rect 11736 23962 11792 23964
rect 11816 23962 11872 23964
rect 11896 23962 11952 23964
rect 11976 23962 12032 23964
rect 11656 23910 11658 23962
rect 11658 23910 11710 23962
rect 11710 23910 11712 23962
rect 11736 23910 11774 23962
rect 11774 23910 11786 23962
rect 11786 23910 11792 23962
rect 11816 23910 11838 23962
rect 11838 23910 11850 23962
rect 11850 23910 11872 23962
rect 11896 23910 11902 23962
rect 11902 23910 11914 23962
rect 11914 23910 11952 23962
rect 11976 23910 11978 23962
rect 11978 23910 12030 23962
rect 12030 23910 12032 23962
rect 11656 23908 11712 23910
rect 11736 23908 11792 23910
rect 11816 23908 11872 23910
rect 11896 23908 11952 23910
rect 11976 23908 12032 23910
rect 11656 22874 11712 22876
rect 11736 22874 11792 22876
rect 11816 22874 11872 22876
rect 11896 22874 11952 22876
rect 11976 22874 12032 22876
rect 11656 22822 11658 22874
rect 11658 22822 11710 22874
rect 11710 22822 11712 22874
rect 11736 22822 11774 22874
rect 11774 22822 11786 22874
rect 11786 22822 11792 22874
rect 11816 22822 11838 22874
rect 11838 22822 11850 22874
rect 11850 22822 11872 22874
rect 11896 22822 11902 22874
rect 11902 22822 11914 22874
rect 11914 22822 11952 22874
rect 11976 22822 11978 22874
rect 11978 22822 12030 22874
rect 12030 22822 12032 22874
rect 11656 22820 11712 22822
rect 11736 22820 11792 22822
rect 11816 22820 11872 22822
rect 11896 22820 11952 22822
rect 11976 22820 12032 22822
rect 10916 22330 10972 22332
rect 10996 22330 11052 22332
rect 11076 22330 11132 22332
rect 11156 22330 11212 22332
rect 11236 22330 11292 22332
rect 10916 22278 10918 22330
rect 10918 22278 10970 22330
rect 10970 22278 10972 22330
rect 10996 22278 11034 22330
rect 11034 22278 11046 22330
rect 11046 22278 11052 22330
rect 11076 22278 11098 22330
rect 11098 22278 11110 22330
rect 11110 22278 11132 22330
rect 11156 22278 11162 22330
rect 11162 22278 11174 22330
rect 11174 22278 11212 22330
rect 11236 22278 11238 22330
rect 11238 22278 11290 22330
rect 11290 22278 11292 22330
rect 10916 22276 10972 22278
rect 10996 22276 11052 22278
rect 11076 22276 11132 22278
rect 11156 22276 11212 22278
rect 11236 22276 11292 22278
rect 11656 21786 11712 21788
rect 11736 21786 11792 21788
rect 11816 21786 11872 21788
rect 11896 21786 11952 21788
rect 11976 21786 12032 21788
rect 11656 21734 11658 21786
rect 11658 21734 11710 21786
rect 11710 21734 11712 21786
rect 11736 21734 11774 21786
rect 11774 21734 11786 21786
rect 11786 21734 11792 21786
rect 11816 21734 11838 21786
rect 11838 21734 11850 21786
rect 11850 21734 11872 21786
rect 11896 21734 11902 21786
rect 11902 21734 11914 21786
rect 11914 21734 11952 21786
rect 11976 21734 11978 21786
rect 11978 21734 12030 21786
rect 12030 21734 12032 21786
rect 11656 21732 11712 21734
rect 11736 21732 11792 21734
rect 11816 21732 11872 21734
rect 11896 21732 11952 21734
rect 11976 21732 12032 21734
rect 10916 21242 10972 21244
rect 10996 21242 11052 21244
rect 11076 21242 11132 21244
rect 11156 21242 11212 21244
rect 11236 21242 11292 21244
rect 10916 21190 10918 21242
rect 10918 21190 10970 21242
rect 10970 21190 10972 21242
rect 10996 21190 11034 21242
rect 11034 21190 11046 21242
rect 11046 21190 11052 21242
rect 11076 21190 11098 21242
rect 11098 21190 11110 21242
rect 11110 21190 11132 21242
rect 11156 21190 11162 21242
rect 11162 21190 11174 21242
rect 11174 21190 11212 21242
rect 11236 21190 11238 21242
rect 11238 21190 11290 21242
rect 11290 21190 11292 21242
rect 10916 21188 10972 21190
rect 10996 21188 11052 21190
rect 11076 21188 11132 21190
rect 11156 21188 11212 21190
rect 11236 21188 11292 21190
rect 11656 20698 11712 20700
rect 11736 20698 11792 20700
rect 11816 20698 11872 20700
rect 11896 20698 11952 20700
rect 11976 20698 12032 20700
rect 11656 20646 11658 20698
rect 11658 20646 11710 20698
rect 11710 20646 11712 20698
rect 11736 20646 11774 20698
rect 11774 20646 11786 20698
rect 11786 20646 11792 20698
rect 11816 20646 11838 20698
rect 11838 20646 11850 20698
rect 11850 20646 11872 20698
rect 11896 20646 11902 20698
rect 11902 20646 11914 20698
rect 11914 20646 11952 20698
rect 11976 20646 11978 20698
rect 11978 20646 12030 20698
rect 12030 20646 12032 20698
rect 11656 20644 11712 20646
rect 11736 20644 11792 20646
rect 11816 20644 11872 20646
rect 11896 20644 11952 20646
rect 11976 20644 12032 20646
rect 10916 20154 10972 20156
rect 10996 20154 11052 20156
rect 11076 20154 11132 20156
rect 11156 20154 11212 20156
rect 11236 20154 11292 20156
rect 10916 20102 10918 20154
rect 10918 20102 10970 20154
rect 10970 20102 10972 20154
rect 10996 20102 11034 20154
rect 11034 20102 11046 20154
rect 11046 20102 11052 20154
rect 11076 20102 11098 20154
rect 11098 20102 11110 20154
rect 11110 20102 11132 20154
rect 11156 20102 11162 20154
rect 11162 20102 11174 20154
rect 11174 20102 11212 20154
rect 11236 20102 11238 20154
rect 11238 20102 11290 20154
rect 11290 20102 11292 20154
rect 10916 20100 10972 20102
rect 10996 20100 11052 20102
rect 11076 20100 11132 20102
rect 11156 20100 11212 20102
rect 11236 20100 11292 20102
rect 11656 19610 11712 19612
rect 11736 19610 11792 19612
rect 11816 19610 11872 19612
rect 11896 19610 11952 19612
rect 11976 19610 12032 19612
rect 11656 19558 11658 19610
rect 11658 19558 11710 19610
rect 11710 19558 11712 19610
rect 11736 19558 11774 19610
rect 11774 19558 11786 19610
rect 11786 19558 11792 19610
rect 11816 19558 11838 19610
rect 11838 19558 11850 19610
rect 11850 19558 11872 19610
rect 11896 19558 11902 19610
rect 11902 19558 11914 19610
rect 11914 19558 11952 19610
rect 11976 19558 11978 19610
rect 11978 19558 12030 19610
rect 12030 19558 12032 19610
rect 11656 19556 11712 19558
rect 11736 19556 11792 19558
rect 11816 19556 11872 19558
rect 11896 19556 11952 19558
rect 11976 19556 12032 19558
rect 10916 19066 10972 19068
rect 10996 19066 11052 19068
rect 11076 19066 11132 19068
rect 11156 19066 11212 19068
rect 11236 19066 11292 19068
rect 10916 19014 10918 19066
rect 10918 19014 10970 19066
rect 10970 19014 10972 19066
rect 10996 19014 11034 19066
rect 11034 19014 11046 19066
rect 11046 19014 11052 19066
rect 11076 19014 11098 19066
rect 11098 19014 11110 19066
rect 11110 19014 11132 19066
rect 11156 19014 11162 19066
rect 11162 19014 11174 19066
rect 11174 19014 11212 19066
rect 11236 19014 11238 19066
rect 11238 19014 11290 19066
rect 11290 19014 11292 19066
rect 10916 19012 10972 19014
rect 10996 19012 11052 19014
rect 11076 19012 11132 19014
rect 11156 19012 11212 19014
rect 11236 19012 11292 19014
rect 10916 17978 10972 17980
rect 10996 17978 11052 17980
rect 11076 17978 11132 17980
rect 11156 17978 11212 17980
rect 11236 17978 11292 17980
rect 10916 17926 10918 17978
rect 10918 17926 10970 17978
rect 10970 17926 10972 17978
rect 10996 17926 11034 17978
rect 11034 17926 11046 17978
rect 11046 17926 11052 17978
rect 11076 17926 11098 17978
rect 11098 17926 11110 17978
rect 11110 17926 11132 17978
rect 11156 17926 11162 17978
rect 11162 17926 11174 17978
rect 11174 17926 11212 17978
rect 11236 17926 11238 17978
rect 11238 17926 11290 17978
rect 11290 17926 11292 17978
rect 10916 17924 10972 17926
rect 10996 17924 11052 17926
rect 11076 17924 11132 17926
rect 11156 17924 11212 17926
rect 11236 17924 11292 17926
rect 12898 23044 12954 23080
rect 12898 23024 12900 23044
rect 12900 23024 12952 23044
rect 12952 23024 12954 23044
rect 15656 27226 15712 27228
rect 15736 27226 15792 27228
rect 15816 27226 15872 27228
rect 15896 27226 15952 27228
rect 15976 27226 16032 27228
rect 15656 27174 15658 27226
rect 15658 27174 15710 27226
rect 15710 27174 15712 27226
rect 15736 27174 15774 27226
rect 15774 27174 15786 27226
rect 15786 27174 15792 27226
rect 15816 27174 15838 27226
rect 15838 27174 15850 27226
rect 15850 27174 15872 27226
rect 15896 27174 15902 27226
rect 15902 27174 15914 27226
rect 15914 27174 15952 27226
rect 15976 27174 15978 27226
rect 15978 27174 16030 27226
rect 16030 27174 16032 27226
rect 15656 27172 15712 27174
rect 15736 27172 15792 27174
rect 15816 27172 15872 27174
rect 15896 27172 15952 27174
rect 15976 27172 16032 27174
rect 11656 18522 11712 18524
rect 11736 18522 11792 18524
rect 11816 18522 11872 18524
rect 11896 18522 11952 18524
rect 11976 18522 12032 18524
rect 11656 18470 11658 18522
rect 11658 18470 11710 18522
rect 11710 18470 11712 18522
rect 11736 18470 11774 18522
rect 11774 18470 11786 18522
rect 11786 18470 11792 18522
rect 11816 18470 11838 18522
rect 11838 18470 11850 18522
rect 11850 18470 11872 18522
rect 11896 18470 11902 18522
rect 11902 18470 11914 18522
rect 11914 18470 11952 18522
rect 11976 18470 11978 18522
rect 11978 18470 12030 18522
rect 12030 18470 12032 18522
rect 11656 18468 11712 18470
rect 11736 18468 11792 18470
rect 11816 18468 11872 18470
rect 11896 18468 11952 18470
rect 11976 18468 12032 18470
rect 10506 15444 10508 15464
rect 10508 15444 10560 15464
rect 10560 15444 10562 15464
rect 10506 15408 10562 15444
rect 10916 16890 10972 16892
rect 10996 16890 11052 16892
rect 11076 16890 11132 16892
rect 11156 16890 11212 16892
rect 11236 16890 11292 16892
rect 10916 16838 10918 16890
rect 10918 16838 10970 16890
rect 10970 16838 10972 16890
rect 10996 16838 11034 16890
rect 11034 16838 11046 16890
rect 11046 16838 11052 16890
rect 11076 16838 11098 16890
rect 11098 16838 11110 16890
rect 11110 16838 11132 16890
rect 11156 16838 11162 16890
rect 11162 16838 11174 16890
rect 11174 16838 11212 16890
rect 11236 16838 11238 16890
rect 11238 16838 11290 16890
rect 11290 16838 11292 16890
rect 10916 16836 10972 16838
rect 10996 16836 11052 16838
rect 11076 16836 11132 16838
rect 11156 16836 11212 16838
rect 11236 16836 11292 16838
rect 11656 17434 11712 17436
rect 11736 17434 11792 17436
rect 11816 17434 11872 17436
rect 11896 17434 11952 17436
rect 11976 17434 12032 17436
rect 11656 17382 11658 17434
rect 11658 17382 11710 17434
rect 11710 17382 11712 17434
rect 11736 17382 11774 17434
rect 11774 17382 11786 17434
rect 11786 17382 11792 17434
rect 11816 17382 11838 17434
rect 11838 17382 11850 17434
rect 11850 17382 11872 17434
rect 11896 17382 11902 17434
rect 11902 17382 11914 17434
rect 11914 17382 11952 17434
rect 11976 17382 11978 17434
rect 11978 17382 12030 17434
rect 12030 17382 12032 17434
rect 11656 17380 11712 17382
rect 11736 17380 11792 17382
rect 11816 17380 11872 17382
rect 11896 17380 11952 17382
rect 11976 17380 12032 17382
rect 11656 16346 11712 16348
rect 11736 16346 11792 16348
rect 11816 16346 11872 16348
rect 11896 16346 11952 16348
rect 11976 16346 12032 16348
rect 11656 16294 11658 16346
rect 11658 16294 11710 16346
rect 11710 16294 11712 16346
rect 11736 16294 11774 16346
rect 11774 16294 11786 16346
rect 11786 16294 11792 16346
rect 11816 16294 11838 16346
rect 11838 16294 11850 16346
rect 11850 16294 11872 16346
rect 11896 16294 11902 16346
rect 11902 16294 11914 16346
rect 11914 16294 11952 16346
rect 11976 16294 11978 16346
rect 11978 16294 12030 16346
rect 12030 16294 12032 16346
rect 11656 16292 11712 16294
rect 11736 16292 11792 16294
rect 11816 16292 11872 16294
rect 11896 16292 11952 16294
rect 11976 16292 12032 16294
rect 10874 15988 10876 16008
rect 10876 15988 10928 16008
rect 10928 15988 10930 16008
rect 10874 15952 10930 15988
rect 10916 15802 10972 15804
rect 10996 15802 11052 15804
rect 11076 15802 11132 15804
rect 11156 15802 11212 15804
rect 11236 15802 11292 15804
rect 10916 15750 10918 15802
rect 10918 15750 10970 15802
rect 10970 15750 10972 15802
rect 10996 15750 11034 15802
rect 11034 15750 11046 15802
rect 11046 15750 11052 15802
rect 11076 15750 11098 15802
rect 11098 15750 11110 15802
rect 11110 15750 11132 15802
rect 11156 15750 11162 15802
rect 11162 15750 11174 15802
rect 11174 15750 11212 15802
rect 11236 15750 11238 15802
rect 11238 15750 11290 15802
rect 11290 15750 11292 15802
rect 10916 15748 10972 15750
rect 10996 15748 11052 15750
rect 11076 15748 11132 15750
rect 11156 15748 11212 15750
rect 11236 15748 11292 15750
rect 11656 15258 11712 15260
rect 11736 15258 11792 15260
rect 11816 15258 11872 15260
rect 11896 15258 11952 15260
rect 11976 15258 12032 15260
rect 11656 15206 11658 15258
rect 11658 15206 11710 15258
rect 11710 15206 11712 15258
rect 11736 15206 11774 15258
rect 11774 15206 11786 15258
rect 11786 15206 11792 15258
rect 11816 15206 11838 15258
rect 11838 15206 11850 15258
rect 11850 15206 11872 15258
rect 11896 15206 11902 15258
rect 11902 15206 11914 15258
rect 11914 15206 11952 15258
rect 11976 15206 11978 15258
rect 11978 15206 12030 15258
rect 12030 15206 12032 15258
rect 11656 15204 11712 15206
rect 11736 15204 11792 15206
rect 11816 15204 11872 15206
rect 11896 15204 11952 15206
rect 11976 15204 12032 15206
rect 11058 15156 11114 15192
rect 11058 15136 11060 15156
rect 11060 15136 11112 15156
rect 11112 15136 11114 15156
rect 10916 14714 10972 14716
rect 10996 14714 11052 14716
rect 11076 14714 11132 14716
rect 11156 14714 11212 14716
rect 11236 14714 11292 14716
rect 10916 14662 10918 14714
rect 10918 14662 10970 14714
rect 10970 14662 10972 14714
rect 10996 14662 11034 14714
rect 11034 14662 11046 14714
rect 11046 14662 11052 14714
rect 11076 14662 11098 14714
rect 11098 14662 11110 14714
rect 11110 14662 11132 14714
rect 11156 14662 11162 14714
rect 11162 14662 11174 14714
rect 11174 14662 11212 14714
rect 11236 14662 11238 14714
rect 11238 14662 11290 14714
rect 11290 14662 11292 14714
rect 10916 14660 10972 14662
rect 10996 14660 11052 14662
rect 11076 14660 11132 14662
rect 11156 14660 11212 14662
rect 11236 14660 11292 14662
rect 11656 14170 11712 14172
rect 11736 14170 11792 14172
rect 11816 14170 11872 14172
rect 11896 14170 11952 14172
rect 11976 14170 12032 14172
rect 11656 14118 11658 14170
rect 11658 14118 11710 14170
rect 11710 14118 11712 14170
rect 11736 14118 11774 14170
rect 11774 14118 11786 14170
rect 11786 14118 11792 14170
rect 11816 14118 11838 14170
rect 11838 14118 11850 14170
rect 11850 14118 11872 14170
rect 11896 14118 11902 14170
rect 11902 14118 11914 14170
rect 11914 14118 11952 14170
rect 11976 14118 11978 14170
rect 11978 14118 12030 14170
rect 12030 14118 12032 14170
rect 11656 14116 11712 14118
rect 11736 14116 11792 14118
rect 11816 14116 11872 14118
rect 11896 14116 11952 14118
rect 11976 14116 12032 14118
rect 10046 10784 10048 10804
rect 10048 10784 10100 10804
rect 10100 10784 10102 10804
rect 7656 5466 7712 5468
rect 7736 5466 7792 5468
rect 7816 5466 7872 5468
rect 7896 5466 7952 5468
rect 7976 5466 8032 5468
rect 7656 5414 7658 5466
rect 7658 5414 7710 5466
rect 7710 5414 7712 5466
rect 7736 5414 7774 5466
rect 7774 5414 7786 5466
rect 7786 5414 7792 5466
rect 7816 5414 7838 5466
rect 7838 5414 7850 5466
rect 7850 5414 7872 5466
rect 7896 5414 7902 5466
rect 7902 5414 7914 5466
rect 7914 5414 7952 5466
rect 7976 5414 7978 5466
rect 7978 5414 8030 5466
rect 8030 5414 8032 5466
rect 7656 5412 7712 5414
rect 7736 5412 7792 5414
rect 7816 5412 7872 5414
rect 7896 5412 7952 5414
rect 7976 5412 8032 5414
rect 7656 4378 7712 4380
rect 7736 4378 7792 4380
rect 7816 4378 7872 4380
rect 7896 4378 7952 4380
rect 7976 4378 8032 4380
rect 7656 4326 7658 4378
rect 7658 4326 7710 4378
rect 7710 4326 7712 4378
rect 7736 4326 7774 4378
rect 7774 4326 7786 4378
rect 7786 4326 7792 4378
rect 7816 4326 7838 4378
rect 7838 4326 7850 4378
rect 7850 4326 7872 4378
rect 7896 4326 7902 4378
rect 7902 4326 7914 4378
rect 7914 4326 7952 4378
rect 7976 4326 7978 4378
rect 7978 4326 8030 4378
rect 8030 4326 8032 4378
rect 7656 4324 7712 4326
rect 7736 4324 7792 4326
rect 7816 4324 7872 4326
rect 7896 4324 7952 4326
rect 7976 4324 8032 4326
rect 7656 3290 7712 3292
rect 7736 3290 7792 3292
rect 7816 3290 7872 3292
rect 7896 3290 7952 3292
rect 7976 3290 8032 3292
rect 7656 3238 7658 3290
rect 7658 3238 7710 3290
rect 7710 3238 7712 3290
rect 7736 3238 7774 3290
rect 7774 3238 7786 3290
rect 7786 3238 7792 3290
rect 7816 3238 7838 3290
rect 7838 3238 7850 3290
rect 7850 3238 7872 3290
rect 7896 3238 7902 3290
rect 7902 3238 7914 3290
rect 7914 3238 7952 3290
rect 7976 3238 7978 3290
rect 7978 3238 8030 3290
rect 8030 3238 8032 3290
rect 7656 3236 7712 3238
rect 7736 3236 7792 3238
rect 7816 3236 7872 3238
rect 7896 3236 7952 3238
rect 7976 3236 8032 3238
rect 10916 13626 10972 13628
rect 10996 13626 11052 13628
rect 11076 13626 11132 13628
rect 11156 13626 11212 13628
rect 11236 13626 11292 13628
rect 10916 13574 10918 13626
rect 10918 13574 10970 13626
rect 10970 13574 10972 13626
rect 10996 13574 11034 13626
rect 11034 13574 11046 13626
rect 11046 13574 11052 13626
rect 11076 13574 11098 13626
rect 11098 13574 11110 13626
rect 11110 13574 11132 13626
rect 11156 13574 11162 13626
rect 11162 13574 11174 13626
rect 11174 13574 11212 13626
rect 11236 13574 11238 13626
rect 11238 13574 11290 13626
rect 11290 13574 11292 13626
rect 10916 13572 10972 13574
rect 10996 13572 11052 13574
rect 11076 13572 11132 13574
rect 11156 13572 11212 13574
rect 11236 13572 11292 13574
rect 10916 12538 10972 12540
rect 10996 12538 11052 12540
rect 11076 12538 11132 12540
rect 11156 12538 11212 12540
rect 11236 12538 11292 12540
rect 10916 12486 10918 12538
rect 10918 12486 10970 12538
rect 10970 12486 10972 12538
rect 10996 12486 11034 12538
rect 11034 12486 11046 12538
rect 11046 12486 11052 12538
rect 11076 12486 11098 12538
rect 11098 12486 11110 12538
rect 11110 12486 11132 12538
rect 11156 12486 11162 12538
rect 11162 12486 11174 12538
rect 11174 12486 11212 12538
rect 11236 12486 11238 12538
rect 11238 12486 11290 12538
rect 11290 12486 11292 12538
rect 10916 12484 10972 12486
rect 10996 12484 11052 12486
rect 11076 12484 11132 12486
rect 11156 12484 11212 12486
rect 11236 12484 11292 12486
rect 10916 11450 10972 11452
rect 10996 11450 11052 11452
rect 11076 11450 11132 11452
rect 11156 11450 11212 11452
rect 11236 11450 11292 11452
rect 10916 11398 10918 11450
rect 10918 11398 10970 11450
rect 10970 11398 10972 11450
rect 10996 11398 11034 11450
rect 11034 11398 11046 11450
rect 11046 11398 11052 11450
rect 11076 11398 11098 11450
rect 11098 11398 11110 11450
rect 11110 11398 11132 11450
rect 11156 11398 11162 11450
rect 11162 11398 11174 11450
rect 11174 11398 11212 11450
rect 11236 11398 11238 11450
rect 11238 11398 11290 11450
rect 11290 11398 11292 11450
rect 10916 11396 10972 11398
rect 10996 11396 11052 11398
rect 11076 11396 11132 11398
rect 11156 11396 11212 11398
rect 11236 11396 11292 11398
rect 10916 10362 10972 10364
rect 10996 10362 11052 10364
rect 11076 10362 11132 10364
rect 11156 10362 11212 10364
rect 11236 10362 11292 10364
rect 10916 10310 10918 10362
rect 10918 10310 10970 10362
rect 10970 10310 10972 10362
rect 10996 10310 11034 10362
rect 11034 10310 11046 10362
rect 11046 10310 11052 10362
rect 11076 10310 11098 10362
rect 11098 10310 11110 10362
rect 11110 10310 11132 10362
rect 11156 10310 11162 10362
rect 11162 10310 11174 10362
rect 11174 10310 11212 10362
rect 11236 10310 11238 10362
rect 11238 10310 11290 10362
rect 11290 10310 11292 10362
rect 10916 10308 10972 10310
rect 10996 10308 11052 10310
rect 11076 10308 11132 10310
rect 11156 10308 11212 10310
rect 11236 10308 11292 10310
rect 11656 13082 11712 13084
rect 11736 13082 11792 13084
rect 11816 13082 11872 13084
rect 11896 13082 11952 13084
rect 11976 13082 12032 13084
rect 11656 13030 11658 13082
rect 11658 13030 11710 13082
rect 11710 13030 11712 13082
rect 11736 13030 11774 13082
rect 11774 13030 11786 13082
rect 11786 13030 11792 13082
rect 11816 13030 11838 13082
rect 11838 13030 11850 13082
rect 11850 13030 11872 13082
rect 11896 13030 11902 13082
rect 11902 13030 11914 13082
rect 11914 13030 11952 13082
rect 11976 13030 11978 13082
rect 11978 13030 12030 13082
rect 12030 13030 12032 13082
rect 11656 13028 11712 13030
rect 11736 13028 11792 13030
rect 11816 13028 11872 13030
rect 11896 13028 11952 13030
rect 11976 13028 12032 13030
rect 11656 11994 11712 11996
rect 11736 11994 11792 11996
rect 11816 11994 11872 11996
rect 11896 11994 11952 11996
rect 11976 11994 12032 11996
rect 11656 11942 11658 11994
rect 11658 11942 11710 11994
rect 11710 11942 11712 11994
rect 11736 11942 11774 11994
rect 11774 11942 11786 11994
rect 11786 11942 11792 11994
rect 11816 11942 11838 11994
rect 11838 11942 11850 11994
rect 11850 11942 11872 11994
rect 11896 11942 11902 11994
rect 11902 11942 11914 11994
rect 11914 11942 11952 11994
rect 11976 11942 11978 11994
rect 11978 11942 12030 11994
rect 12030 11942 12032 11994
rect 11656 11940 11712 11942
rect 11736 11940 11792 11942
rect 11816 11940 11872 11942
rect 11896 11940 11952 11942
rect 11976 11940 12032 11942
rect 11656 10906 11712 10908
rect 11736 10906 11792 10908
rect 11816 10906 11872 10908
rect 11896 10906 11952 10908
rect 11976 10906 12032 10908
rect 11656 10854 11658 10906
rect 11658 10854 11710 10906
rect 11710 10854 11712 10906
rect 11736 10854 11774 10906
rect 11774 10854 11786 10906
rect 11786 10854 11792 10906
rect 11816 10854 11838 10906
rect 11838 10854 11850 10906
rect 11850 10854 11872 10906
rect 11896 10854 11902 10906
rect 11902 10854 11914 10906
rect 11914 10854 11952 10906
rect 11976 10854 11978 10906
rect 11978 10854 12030 10906
rect 12030 10854 12032 10906
rect 11656 10852 11712 10854
rect 11736 10852 11792 10854
rect 11816 10852 11872 10854
rect 11896 10852 11952 10854
rect 11976 10852 12032 10854
rect 10598 8472 10654 8528
rect 10916 9274 10972 9276
rect 10996 9274 11052 9276
rect 11076 9274 11132 9276
rect 11156 9274 11212 9276
rect 11236 9274 11292 9276
rect 10916 9222 10918 9274
rect 10918 9222 10970 9274
rect 10970 9222 10972 9274
rect 10996 9222 11034 9274
rect 11034 9222 11046 9274
rect 11046 9222 11052 9274
rect 11076 9222 11098 9274
rect 11098 9222 11110 9274
rect 11110 9222 11132 9274
rect 11156 9222 11162 9274
rect 11162 9222 11174 9274
rect 11174 9222 11212 9274
rect 11236 9222 11238 9274
rect 11238 9222 11290 9274
rect 11290 9222 11292 9274
rect 10916 9220 10972 9222
rect 10996 9220 11052 9222
rect 11076 9220 11132 9222
rect 11156 9220 11212 9222
rect 11236 9220 11292 9222
rect 10916 8186 10972 8188
rect 10996 8186 11052 8188
rect 11076 8186 11132 8188
rect 11156 8186 11212 8188
rect 11236 8186 11292 8188
rect 10916 8134 10918 8186
rect 10918 8134 10970 8186
rect 10970 8134 10972 8186
rect 10996 8134 11034 8186
rect 11034 8134 11046 8186
rect 11046 8134 11052 8186
rect 11076 8134 11098 8186
rect 11098 8134 11110 8186
rect 11110 8134 11132 8186
rect 11156 8134 11162 8186
rect 11162 8134 11174 8186
rect 11174 8134 11212 8186
rect 11236 8134 11238 8186
rect 11238 8134 11290 8186
rect 11290 8134 11292 8186
rect 10916 8132 10972 8134
rect 10996 8132 11052 8134
rect 11076 8132 11132 8134
rect 11156 8132 11212 8134
rect 11236 8132 11292 8134
rect 11656 9818 11712 9820
rect 11736 9818 11792 9820
rect 11816 9818 11872 9820
rect 11896 9818 11952 9820
rect 11976 9818 12032 9820
rect 11656 9766 11658 9818
rect 11658 9766 11710 9818
rect 11710 9766 11712 9818
rect 11736 9766 11774 9818
rect 11774 9766 11786 9818
rect 11786 9766 11792 9818
rect 11816 9766 11838 9818
rect 11838 9766 11850 9818
rect 11850 9766 11872 9818
rect 11896 9766 11902 9818
rect 11902 9766 11914 9818
rect 11914 9766 11952 9818
rect 11976 9766 11978 9818
rect 11978 9766 12030 9818
rect 12030 9766 12032 9818
rect 11656 9764 11712 9766
rect 11736 9764 11792 9766
rect 11816 9764 11872 9766
rect 11896 9764 11952 9766
rect 11976 9764 12032 9766
rect 11656 8730 11712 8732
rect 11736 8730 11792 8732
rect 11816 8730 11872 8732
rect 11896 8730 11952 8732
rect 11976 8730 12032 8732
rect 11656 8678 11658 8730
rect 11658 8678 11710 8730
rect 11710 8678 11712 8730
rect 11736 8678 11774 8730
rect 11774 8678 11786 8730
rect 11786 8678 11792 8730
rect 11816 8678 11838 8730
rect 11838 8678 11850 8730
rect 11850 8678 11872 8730
rect 11896 8678 11902 8730
rect 11902 8678 11914 8730
rect 11914 8678 11952 8730
rect 11976 8678 11978 8730
rect 11978 8678 12030 8730
rect 12030 8678 12032 8730
rect 11656 8676 11712 8678
rect 11736 8676 11792 8678
rect 11816 8676 11872 8678
rect 11896 8676 11952 8678
rect 11976 8676 12032 8678
rect 12898 17076 12900 17096
rect 12900 17076 12952 17096
rect 12952 17076 12954 17096
rect 12898 17040 12954 17076
rect 14916 26682 14972 26684
rect 14996 26682 15052 26684
rect 15076 26682 15132 26684
rect 15156 26682 15212 26684
rect 15236 26682 15292 26684
rect 14916 26630 14918 26682
rect 14918 26630 14970 26682
rect 14970 26630 14972 26682
rect 14996 26630 15034 26682
rect 15034 26630 15046 26682
rect 15046 26630 15052 26682
rect 15076 26630 15098 26682
rect 15098 26630 15110 26682
rect 15110 26630 15132 26682
rect 15156 26630 15162 26682
rect 15162 26630 15174 26682
rect 15174 26630 15212 26682
rect 15236 26630 15238 26682
rect 15238 26630 15290 26682
rect 15290 26630 15292 26682
rect 14916 26628 14972 26630
rect 14996 26628 15052 26630
rect 15076 26628 15132 26630
rect 15156 26628 15212 26630
rect 15236 26628 15292 26630
rect 15656 26138 15712 26140
rect 15736 26138 15792 26140
rect 15816 26138 15872 26140
rect 15896 26138 15952 26140
rect 15976 26138 16032 26140
rect 15656 26086 15658 26138
rect 15658 26086 15710 26138
rect 15710 26086 15712 26138
rect 15736 26086 15774 26138
rect 15774 26086 15786 26138
rect 15786 26086 15792 26138
rect 15816 26086 15838 26138
rect 15838 26086 15850 26138
rect 15850 26086 15872 26138
rect 15896 26086 15902 26138
rect 15902 26086 15914 26138
rect 15914 26086 15952 26138
rect 15976 26086 15978 26138
rect 15978 26086 16030 26138
rect 16030 26086 16032 26138
rect 15656 26084 15712 26086
rect 15736 26084 15792 26086
rect 15816 26084 15872 26086
rect 15896 26084 15952 26086
rect 15976 26084 16032 26086
rect 14916 25594 14972 25596
rect 14996 25594 15052 25596
rect 15076 25594 15132 25596
rect 15156 25594 15212 25596
rect 15236 25594 15292 25596
rect 14916 25542 14918 25594
rect 14918 25542 14970 25594
rect 14970 25542 14972 25594
rect 14996 25542 15034 25594
rect 15034 25542 15046 25594
rect 15046 25542 15052 25594
rect 15076 25542 15098 25594
rect 15098 25542 15110 25594
rect 15110 25542 15132 25594
rect 15156 25542 15162 25594
rect 15162 25542 15174 25594
rect 15174 25542 15212 25594
rect 15236 25542 15238 25594
rect 15238 25542 15290 25594
rect 15290 25542 15292 25594
rect 14916 25540 14972 25542
rect 14996 25540 15052 25542
rect 15076 25540 15132 25542
rect 15156 25540 15212 25542
rect 15236 25540 15292 25542
rect 15656 25050 15712 25052
rect 15736 25050 15792 25052
rect 15816 25050 15872 25052
rect 15896 25050 15952 25052
rect 15976 25050 16032 25052
rect 15656 24998 15658 25050
rect 15658 24998 15710 25050
rect 15710 24998 15712 25050
rect 15736 24998 15774 25050
rect 15774 24998 15786 25050
rect 15786 24998 15792 25050
rect 15816 24998 15838 25050
rect 15838 24998 15850 25050
rect 15850 24998 15872 25050
rect 15896 24998 15902 25050
rect 15902 24998 15914 25050
rect 15914 24998 15952 25050
rect 15976 24998 15978 25050
rect 15978 24998 16030 25050
rect 16030 24998 16032 25050
rect 15656 24996 15712 24998
rect 15736 24996 15792 24998
rect 15816 24996 15872 24998
rect 15896 24996 15952 24998
rect 15976 24996 16032 24998
rect 14916 24506 14972 24508
rect 14996 24506 15052 24508
rect 15076 24506 15132 24508
rect 15156 24506 15212 24508
rect 15236 24506 15292 24508
rect 14916 24454 14918 24506
rect 14918 24454 14970 24506
rect 14970 24454 14972 24506
rect 14996 24454 15034 24506
rect 15034 24454 15046 24506
rect 15046 24454 15052 24506
rect 15076 24454 15098 24506
rect 15098 24454 15110 24506
rect 15110 24454 15132 24506
rect 15156 24454 15162 24506
rect 15162 24454 15174 24506
rect 15174 24454 15212 24506
rect 15236 24454 15238 24506
rect 15238 24454 15290 24506
rect 15290 24454 15292 24506
rect 14916 24452 14972 24454
rect 14996 24452 15052 24454
rect 15076 24452 15132 24454
rect 15156 24452 15212 24454
rect 15236 24452 15292 24454
rect 15656 23962 15712 23964
rect 15736 23962 15792 23964
rect 15816 23962 15872 23964
rect 15896 23962 15952 23964
rect 15976 23962 16032 23964
rect 15656 23910 15658 23962
rect 15658 23910 15710 23962
rect 15710 23910 15712 23962
rect 15736 23910 15774 23962
rect 15774 23910 15786 23962
rect 15786 23910 15792 23962
rect 15816 23910 15838 23962
rect 15838 23910 15850 23962
rect 15850 23910 15872 23962
rect 15896 23910 15902 23962
rect 15902 23910 15914 23962
rect 15914 23910 15952 23962
rect 15976 23910 15978 23962
rect 15978 23910 16030 23962
rect 16030 23910 16032 23962
rect 15656 23908 15712 23910
rect 15736 23908 15792 23910
rect 15816 23908 15872 23910
rect 15896 23908 15952 23910
rect 15976 23908 16032 23910
rect 14916 23418 14972 23420
rect 14996 23418 15052 23420
rect 15076 23418 15132 23420
rect 15156 23418 15212 23420
rect 15236 23418 15292 23420
rect 14916 23366 14918 23418
rect 14918 23366 14970 23418
rect 14970 23366 14972 23418
rect 14996 23366 15034 23418
rect 15034 23366 15046 23418
rect 15046 23366 15052 23418
rect 15076 23366 15098 23418
rect 15098 23366 15110 23418
rect 15110 23366 15132 23418
rect 15156 23366 15162 23418
rect 15162 23366 15174 23418
rect 15174 23366 15212 23418
rect 15236 23366 15238 23418
rect 15238 23366 15290 23418
rect 15290 23366 15292 23418
rect 14916 23364 14972 23366
rect 14996 23364 15052 23366
rect 15076 23364 15132 23366
rect 15156 23364 15212 23366
rect 15236 23364 15292 23366
rect 13634 16532 13636 16552
rect 13636 16532 13688 16552
rect 13688 16532 13690 16552
rect 13634 16496 13690 16532
rect 13450 14320 13506 14376
rect 11242 7792 11298 7848
rect 10916 7098 10972 7100
rect 10996 7098 11052 7100
rect 11076 7098 11132 7100
rect 11156 7098 11212 7100
rect 11236 7098 11292 7100
rect 10916 7046 10918 7098
rect 10918 7046 10970 7098
rect 10970 7046 10972 7098
rect 10996 7046 11034 7098
rect 11034 7046 11046 7098
rect 11046 7046 11052 7098
rect 11076 7046 11098 7098
rect 11098 7046 11110 7098
rect 11110 7046 11132 7098
rect 11156 7046 11162 7098
rect 11162 7046 11174 7098
rect 11174 7046 11212 7098
rect 11236 7046 11238 7098
rect 11238 7046 11290 7098
rect 11290 7046 11292 7098
rect 10916 7044 10972 7046
rect 10996 7044 11052 7046
rect 11076 7044 11132 7046
rect 11156 7044 11212 7046
rect 11236 7044 11292 7046
rect 10916 6010 10972 6012
rect 10996 6010 11052 6012
rect 11076 6010 11132 6012
rect 11156 6010 11212 6012
rect 11236 6010 11292 6012
rect 10916 5958 10918 6010
rect 10918 5958 10970 6010
rect 10970 5958 10972 6010
rect 10996 5958 11034 6010
rect 11034 5958 11046 6010
rect 11046 5958 11052 6010
rect 11076 5958 11098 6010
rect 11098 5958 11110 6010
rect 11110 5958 11132 6010
rect 11156 5958 11162 6010
rect 11162 5958 11174 6010
rect 11174 5958 11212 6010
rect 11236 5958 11238 6010
rect 11238 5958 11290 6010
rect 11290 5958 11292 6010
rect 10916 5956 10972 5958
rect 10996 5956 11052 5958
rect 11076 5956 11132 5958
rect 11156 5956 11212 5958
rect 11236 5956 11292 5958
rect 10916 4922 10972 4924
rect 10996 4922 11052 4924
rect 11076 4922 11132 4924
rect 11156 4922 11212 4924
rect 11236 4922 11292 4924
rect 10916 4870 10918 4922
rect 10918 4870 10970 4922
rect 10970 4870 10972 4922
rect 10996 4870 11034 4922
rect 11034 4870 11046 4922
rect 11046 4870 11052 4922
rect 11076 4870 11098 4922
rect 11098 4870 11110 4922
rect 11110 4870 11132 4922
rect 11156 4870 11162 4922
rect 11162 4870 11174 4922
rect 11174 4870 11212 4922
rect 11236 4870 11238 4922
rect 11238 4870 11290 4922
rect 11290 4870 11292 4922
rect 10916 4868 10972 4870
rect 10996 4868 11052 4870
rect 11076 4868 11132 4870
rect 11156 4868 11212 4870
rect 11236 4868 11292 4870
rect 11656 7642 11712 7644
rect 11736 7642 11792 7644
rect 11816 7642 11872 7644
rect 11896 7642 11952 7644
rect 11976 7642 12032 7644
rect 11656 7590 11658 7642
rect 11658 7590 11710 7642
rect 11710 7590 11712 7642
rect 11736 7590 11774 7642
rect 11774 7590 11786 7642
rect 11786 7590 11792 7642
rect 11816 7590 11838 7642
rect 11838 7590 11850 7642
rect 11850 7590 11872 7642
rect 11896 7590 11902 7642
rect 11902 7590 11914 7642
rect 11914 7590 11952 7642
rect 11976 7590 11978 7642
rect 11978 7590 12030 7642
rect 12030 7590 12032 7642
rect 11656 7588 11712 7590
rect 11736 7588 11792 7590
rect 11816 7588 11872 7590
rect 11896 7588 11952 7590
rect 11976 7588 12032 7590
rect 11656 6554 11712 6556
rect 11736 6554 11792 6556
rect 11816 6554 11872 6556
rect 11896 6554 11952 6556
rect 11976 6554 12032 6556
rect 11656 6502 11658 6554
rect 11658 6502 11710 6554
rect 11710 6502 11712 6554
rect 11736 6502 11774 6554
rect 11774 6502 11786 6554
rect 11786 6502 11792 6554
rect 11816 6502 11838 6554
rect 11838 6502 11850 6554
rect 11850 6502 11872 6554
rect 11896 6502 11902 6554
rect 11902 6502 11914 6554
rect 11914 6502 11952 6554
rect 11976 6502 11978 6554
rect 11978 6502 12030 6554
rect 12030 6502 12032 6554
rect 11656 6500 11712 6502
rect 11736 6500 11792 6502
rect 11816 6500 11872 6502
rect 11896 6500 11952 6502
rect 11976 6500 12032 6502
rect 14002 15036 14004 15056
rect 14004 15036 14056 15056
rect 14056 15036 14058 15056
rect 14002 15000 14058 15036
rect 14916 22330 14972 22332
rect 14996 22330 15052 22332
rect 15076 22330 15132 22332
rect 15156 22330 15212 22332
rect 15236 22330 15292 22332
rect 14916 22278 14918 22330
rect 14918 22278 14970 22330
rect 14970 22278 14972 22330
rect 14996 22278 15034 22330
rect 15034 22278 15046 22330
rect 15046 22278 15052 22330
rect 15076 22278 15098 22330
rect 15098 22278 15110 22330
rect 15110 22278 15132 22330
rect 15156 22278 15162 22330
rect 15162 22278 15174 22330
rect 15174 22278 15212 22330
rect 15236 22278 15238 22330
rect 15238 22278 15290 22330
rect 15290 22278 15292 22330
rect 14916 22276 14972 22278
rect 14996 22276 15052 22278
rect 15076 22276 15132 22278
rect 15156 22276 15212 22278
rect 15236 22276 15292 22278
rect 15656 22874 15712 22876
rect 15736 22874 15792 22876
rect 15816 22874 15872 22876
rect 15896 22874 15952 22876
rect 15976 22874 16032 22876
rect 15656 22822 15658 22874
rect 15658 22822 15710 22874
rect 15710 22822 15712 22874
rect 15736 22822 15774 22874
rect 15774 22822 15786 22874
rect 15786 22822 15792 22874
rect 15816 22822 15838 22874
rect 15838 22822 15850 22874
rect 15850 22822 15872 22874
rect 15896 22822 15902 22874
rect 15902 22822 15914 22874
rect 15914 22822 15952 22874
rect 15976 22822 15978 22874
rect 15978 22822 16030 22874
rect 16030 22822 16032 22874
rect 15656 22820 15712 22822
rect 15736 22820 15792 22822
rect 15816 22820 15872 22822
rect 15896 22820 15952 22822
rect 15976 22820 16032 22822
rect 14916 21242 14972 21244
rect 14996 21242 15052 21244
rect 15076 21242 15132 21244
rect 15156 21242 15212 21244
rect 15236 21242 15292 21244
rect 14916 21190 14918 21242
rect 14918 21190 14970 21242
rect 14970 21190 14972 21242
rect 14996 21190 15034 21242
rect 15034 21190 15046 21242
rect 15046 21190 15052 21242
rect 15076 21190 15098 21242
rect 15098 21190 15110 21242
rect 15110 21190 15132 21242
rect 15156 21190 15162 21242
rect 15162 21190 15174 21242
rect 15174 21190 15212 21242
rect 15236 21190 15238 21242
rect 15238 21190 15290 21242
rect 15290 21190 15292 21242
rect 14916 21188 14972 21190
rect 14996 21188 15052 21190
rect 15076 21188 15132 21190
rect 15156 21188 15212 21190
rect 15236 21188 15292 21190
rect 15656 21786 15712 21788
rect 15736 21786 15792 21788
rect 15816 21786 15872 21788
rect 15896 21786 15952 21788
rect 15976 21786 16032 21788
rect 15656 21734 15658 21786
rect 15658 21734 15710 21786
rect 15710 21734 15712 21786
rect 15736 21734 15774 21786
rect 15774 21734 15786 21786
rect 15786 21734 15792 21786
rect 15816 21734 15838 21786
rect 15838 21734 15850 21786
rect 15850 21734 15872 21786
rect 15896 21734 15902 21786
rect 15902 21734 15914 21786
rect 15914 21734 15952 21786
rect 15976 21734 15978 21786
rect 15978 21734 16030 21786
rect 16030 21734 16032 21786
rect 15656 21732 15712 21734
rect 15736 21732 15792 21734
rect 15816 21732 15872 21734
rect 15896 21732 15952 21734
rect 15976 21732 16032 21734
rect 15474 20304 15530 20360
rect 14916 20154 14972 20156
rect 14996 20154 15052 20156
rect 15076 20154 15132 20156
rect 15156 20154 15212 20156
rect 15236 20154 15292 20156
rect 14916 20102 14918 20154
rect 14918 20102 14970 20154
rect 14970 20102 14972 20154
rect 14996 20102 15034 20154
rect 15034 20102 15046 20154
rect 15046 20102 15052 20154
rect 15076 20102 15098 20154
rect 15098 20102 15110 20154
rect 15110 20102 15132 20154
rect 15156 20102 15162 20154
rect 15162 20102 15174 20154
rect 15174 20102 15212 20154
rect 15236 20102 15238 20154
rect 15238 20102 15290 20154
rect 15290 20102 15292 20154
rect 14916 20100 14972 20102
rect 14996 20100 15052 20102
rect 15076 20100 15132 20102
rect 15156 20100 15212 20102
rect 15236 20100 15292 20102
rect 14916 19066 14972 19068
rect 14996 19066 15052 19068
rect 15076 19066 15132 19068
rect 15156 19066 15212 19068
rect 15236 19066 15292 19068
rect 14916 19014 14918 19066
rect 14918 19014 14970 19066
rect 14970 19014 14972 19066
rect 14996 19014 15034 19066
rect 15034 19014 15046 19066
rect 15046 19014 15052 19066
rect 15076 19014 15098 19066
rect 15098 19014 15110 19066
rect 15110 19014 15132 19066
rect 15156 19014 15162 19066
rect 15162 19014 15174 19066
rect 15174 19014 15212 19066
rect 15236 19014 15238 19066
rect 15238 19014 15290 19066
rect 15290 19014 15292 19066
rect 14916 19012 14972 19014
rect 14996 19012 15052 19014
rect 15076 19012 15132 19014
rect 15156 19012 15212 19014
rect 15236 19012 15292 19014
rect 14916 17978 14972 17980
rect 14996 17978 15052 17980
rect 15076 17978 15132 17980
rect 15156 17978 15212 17980
rect 15236 17978 15292 17980
rect 14916 17926 14918 17978
rect 14918 17926 14970 17978
rect 14970 17926 14972 17978
rect 14996 17926 15034 17978
rect 15034 17926 15046 17978
rect 15046 17926 15052 17978
rect 15076 17926 15098 17978
rect 15098 17926 15110 17978
rect 15110 17926 15132 17978
rect 15156 17926 15162 17978
rect 15162 17926 15174 17978
rect 15174 17926 15212 17978
rect 15236 17926 15238 17978
rect 15238 17926 15290 17978
rect 15290 17926 15292 17978
rect 14916 17924 14972 17926
rect 14996 17924 15052 17926
rect 15076 17924 15132 17926
rect 15156 17924 15212 17926
rect 15236 17924 15292 17926
rect 14916 16890 14972 16892
rect 14996 16890 15052 16892
rect 15076 16890 15132 16892
rect 15156 16890 15212 16892
rect 15236 16890 15292 16892
rect 14916 16838 14918 16890
rect 14918 16838 14970 16890
rect 14970 16838 14972 16890
rect 14996 16838 15034 16890
rect 15034 16838 15046 16890
rect 15046 16838 15052 16890
rect 15076 16838 15098 16890
rect 15098 16838 15110 16890
rect 15110 16838 15132 16890
rect 15156 16838 15162 16890
rect 15162 16838 15174 16890
rect 15174 16838 15212 16890
rect 15236 16838 15238 16890
rect 15238 16838 15290 16890
rect 15290 16838 15292 16890
rect 14916 16836 14972 16838
rect 14996 16836 15052 16838
rect 15076 16836 15132 16838
rect 15156 16836 15212 16838
rect 15236 16836 15292 16838
rect 14916 15802 14972 15804
rect 14996 15802 15052 15804
rect 15076 15802 15132 15804
rect 15156 15802 15212 15804
rect 15236 15802 15292 15804
rect 14916 15750 14918 15802
rect 14918 15750 14970 15802
rect 14970 15750 14972 15802
rect 14996 15750 15034 15802
rect 15034 15750 15046 15802
rect 15046 15750 15052 15802
rect 15076 15750 15098 15802
rect 15098 15750 15110 15802
rect 15110 15750 15132 15802
rect 15156 15750 15162 15802
rect 15162 15750 15174 15802
rect 15174 15750 15212 15802
rect 15236 15750 15238 15802
rect 15238 15750 15290 15802
rect 15290 15750 15292 15802
rect 14916 15748 14972 15750
rect 14996 15748 15052 15750
rect 15076 15748 15132 15750
rect 15156 15748 15212 15750
rect 15236 15748 15292 15750
rect 14916 14714 14972 14716
rect 14996 14714 15052 14716
rect 15076 14714 15132 14716
rect 15156 14714 15212 14716
rect 15236 14714 15292 14716
rect 14916 14662 14918 14714
rect 14918 14662 14970 14714
rect 14970 14662 14972 14714
rect 14996 14662 15034 14714
rect 15034 14662 15046 14714
rect 15046 14662 15052 14714
rect 15076 14662 15098 14714
rect 15098 14662 15110 14714
rect 15110 14662 15132 14714
rect 15156 14662 15162 14714
rect 15162 14662 15174 14714
rect 15174 14662 15212 14714
rect 15236 14662 15238 14714
rect 15238 14662 15290 14714
rect 15290 14662 15292 14714
rect 14916 14660 14972 14662
rect 14996 14660 15052 14662
rect 15076 14660 15132 14662
rect 15156 14660 15212 14662
rect 15236 14660 15292 14662
rect 14830 14456 14886 14512
rect 15656 20698 15712 20700
rect 15736 20698 15792 20700
rect 15816 20698 15872 20700
rect 15896 20698 15952 20700
rect 15976 20698 16032 20700
rect 15656 20646 15658 20698
rect 15658 20646 15710 20698
rect 15710 20646 15712 20698
rect 15736 20646 15774 20698
rect 15774 20646 15786 20698
rect 15786 20646 15792 20698
rect 15816 20646 15838 20698
rect 15838 20646 15850 20698
rect 15850 20646 15872 20698
rect 15896 20646 15902 20698
rect 15902 20646 15914 20698
rect 15914 20646 15952 20698
rect 15976 20646 15978 20698
rect 15978 20646 16030 20698
rect 16030 20646 16032 20698
rect 15656 20644 15712 20646
rect 15736 20644 15792 20646
rect 15816 20644 15872 20646
rect 15896 20644 15952 20646
rect 15976 20644 16032 20646
rect 15656 19610 15712 19612
rect 15736 19610 15792 19612
rect 15816 19610 15872 19612
rect 15896 19610 15952 19612
rect 15976 19610 16032 19612
rect 15656 19558 15658 19610
rect 15658 19558 15710 19610
rect 15710 19558 15712 19610
rect 15736 19558 15774 19610
rect 15774 19558 15786 19610
rect 15786 19558 15792 19610
rect 15816 19558 15838 19610
rect 15838 19558 15850 19610
rect 15850 19558 15872 19610
rect 15896 19558 15902 19610
rect 15902 19558 15914 19610
rect 15914 19558 15952 19610
rect 15976 19558 15978 19610
rect 15978 19558 16030 19610
rect 16030 19558 16032 19610
rect 15656 19556 15712 19558
rect 15736 19556 15792 19558
rect 15816 19556 15872 19558
rect 15896 19556 15952 19558
rect 15976 19556 16032 19558
rect 15656 18522 15712 18524
rect 15736 18522 15792 18524
rect 15816 18522 15872 18524
rect 15896 18522 15952 18524
rect 15976 18522 16032 18524
rect 15656 18470 15658 18522
rect 15658 18470 15710 18522
rect 15710 18470 15712 18522
rect 15736 18470 15774 18522
rect 15774 18470 15786 18522
rect 15786 18470 15792 18522
rect 15816 18470 15838 18522
rect 15838 18470 15850 18522
rect 15850 18470 15872 18522
rect 15896 18470 15902 18522
rect 15902 18470 15914 18522
rect 15914 18470 15952 18522
rect 15976 18470 15978 18522
rect 15978 18470 16030 18522
rect 16030 18470 16032 18522
rect 15656 18468 15712 18470
rect 15736 18468 15792 18470
rect 15816 18468 15872 18470
rect 15896 18468 15952 18470
rect 15976 18468 16032 18470
rect 15656 17434 15712 17436
rect 15736 17434 15792 17436
rect 15816 17434 15872 17436
rect 15896 17434 15952 17436
rect 15976 17434 16032 17436
rect 15656 17382 15658 17434
rect 15658 17382 15710 17434
rect 15710 17382 15712 17434
rect 15736 17382 15774 17434
rect 15774 17382 15786 17434
rect 15786 17382 15792 17434
rect 15816 17382 15838 17434
rect 15838 17382 15850 17434
rect 15850 17382 15872 17434
rect 15896 17382 15902 17434
rect 15902 17382 15914 17434
rect 15914 17382 15952 17434
rect 15976 17382 15978 17434
rect 15978 17382 16030 17434
rect 16030 17382 16032 17434
rect 15656 17380 15712 17382
rect 15736 17380 15792 17382
rect 15816 17380 15872 17382
rect 15896 17380 15952 17382
rect 15976 17380 16032 17382
rect 15566 16632 15622 16688
rect 15656 16346 15712 16348
rect 15736 16346 15792 16348
rect 15816 16346 15872 16348
rect 15896 16346 15952 16348
rect 15976 16346 16032 16348
rect 15656 16294 15658 16346
rect 15658 16294 15710 16346
rect 15710 16294 15712 16346
rect 15736 16294 15774 16346
rect 15774 16294 15786 16346
rect 15786 16294 15792 16346
rect 15816 16294 15838 16346
rect 15838 16294 15850 16346
rect 15850 16294 15872 16346
rect 15896 16294 15902 16346
rect 15902 16294 15914 16346
rect 15914 16294 15952 16346
rect 15976 16294 15978 16346
rect 15978 16294 16030 16346
rect 16030 16294 16032 16346
rect 15656 16292 15712 16294
rect 15736 16292 15792 16294
rect 15816 16292 15872 16294
rect 15896 16292 15952 16294
rect 15976 16292 16032 16294
rect 14916 13626 14972 13628
rect 14996 13626 15052 13628
rect 15076 13626 15132 13628
rect 15156 13626 15212 13628
rect 15236 13626 15292 13628
rect 14916 13574 14918 13626
rect 14918 13574 14970 13626
rect 14970 13574 14972 13626
rect 14996 13574 15034 13626
rect 15034 13574 15046 13626
rect 15046 13574 15052 13626
rect 15076 13574 15098 13626
rect 15098 13574 15110 13626
rect 15110 13574 15132 13626
rect 15156 13574 15162 13626
rect 15162 13574 15174 13626
rect 15174 13574 15212 13626
rect 15236 13574 15238 13626
rect 15238 13574 15290 13626
rect 15290 13574 15292 13626
rect 14916 13572 14972 13574
rect 14996 13572 15052 13574
rect 15076 13572 15132 13574
rect 15156 13572 15212 13574
rect 15236 13572 15292 13574
rect 14916 12538 14972 12540
rect 14996 12538 15052 12540
rect 15076 12538 15132 12540
rect 15156 12538 15212 12540
rect 15236 12538 15292 12540
rect 14916 12486 14918 12538
rect 14918 12486 14970 12538
rect 14970 12486 14972 12538
rect 14996 12486 15034 12538
rect 15034 12486 15046 12538
rect 15046 12486 15052 12538
rect 15076 12486 15098 12538
rect 15098 12486 15110 12538
rect 15110 12486 15132 12538
rect 15156 12486 15162 12538
rect 15162 12486 15174 12538
rect 15174 12486 15212 12538
rect 15236 12486 15238 12538
rect 15238 12486 15290 12538
rect 15290 12486 15292 12538
rect 14916 12484 14972 12486
rect 14996 12484 15052 12486
rect 15076 12484 15132 12486
rect 15156 12484 15212 12486
rect 15236 12484 15292 12486
rect 14916 11450 14972 11452
rect 14996 11450 15052 11452
rect 15076 11450 15132 11452
rect 15156 11450 15212 11452
rect 15236 11450 15292 11452
rect 14916 11398 14918 11450
rect 14918 11398 14970 11450
rect 14970 11398 14972 11450
rect 14996 11398 15034 11450
rect 15034 11398 15046 11450
rect 15046 11398 15052 11450
rect 15076 11398 15098 11450
rect 15098 11398 15110 11450
rect 15110 11398 15132 11450
rect 15156 11398 15162 11450
rect 15162 11398 15174 11450
rect 15174 11398 15212 11450
rect 15236 11398 15238 11450
rect 15238 11398 15290 11450
rect 15290 11398 15292 11450
rect 14916 11396 14972 11398
rect 14996 11396 15052 11398
rect 15076 11396 15132 11398
rect 15156 11396 15212 11398
rect 15236 11396 15292 11398
rect 14278 10004 14280 10024
rect 14280 10004 14332 10024
rect 14332 10004 14334 10024
rect 14278 9968 14334 10004
rect 14554 8492 14610 8528
rect 14554 8472 14556 8492
rect 14556 8472 14608 8492
rect 14608 8472 14610 8492
rect 11656 5466 11712 5468
rect 11736 5466 11792 5468
rect 11816 5466 11872 5468
rect 11896 5466 11952 5468
rect 11976 5466 12032 5468
rect 11656 5414 11658 5466
rect 11658 5414 11710 5466
rect 11710 5414 11712 5466
rect 11736 5414 11774 5466
rect 11774 5414 11786 5466
rect 11786 5414 11792 5466
rect 11816 5414 11838 5466
rect 11838 5414 11850 5466
rect 11850 5414 11872 5466
rect 11896 5414 11902 5466
rect 11902 5414 11914 5466
rect 11914 5414 11952 5466
rect 11976 5414 11978 5466
rect 11978 5414 12030 5466
rect 12030 5414 12032 5466
rect 11656 5412 11712 5414
rect 11736 5412 11792 5414
rect 11816 5412 11872 5414
rect 11896 5412 11952 5414
rect 11976 5412 12032 5414
rect 11656 4378 11712 4380
rect 11736 4378 11792 4380
rect 11816 4378 11872 4380
rect 11896 4378 11952 4380
rect 11976 4378 12032 4380
rect 11656 4326 11658 4378
rect 11658 4326 11710 4378
rect 11710 4326 11712 4378
rect 11736 4326 11774 4378
rect 11774 4326 11786 4378
rect 11786 4326 11792 4378
rect 11816 4326 11838 4378
rect 11838 4326 11850 4378
rect 11850 4326 11872 4378
rect 11896 4326 11902 4378
rect 11902 4326 11914 4378
rect 11914 4326 11952 4378
rect 11976 4326 11978 4378
rect 11978 4326 12030 4378
rect 12030 4326 12032 4378
rect 11656 4324 11712 4326
rect 11736 4324 11792 4326
rect 11816 4324 11872 4326
rect 11896 4324 11952 4326
rect 11976 4324 12032 4326
rect 10916 3834 10972 3836
rect 10996 3834 11052 3836
rect 11076 3834 11132 3836
rect 11156 3834 11212 3836
rect 11236 3834 11292 3836
rect 10916 3782 10918 3834
rect 10918 3782 10970 3834
rect 10970 3782 10972 3834
rect 10996 3782 11034 3834
rect 11034 3782 11046 3834
rect 11046 3782 11052 3834
rect 11076 3782 11098 3834
rect 11098 3782 11110 3834
rect 11110 3782 11132 3834
rect 11156 3782 11162 3834
rect 11162 3782 11174 3834
rect 11174 3782 11212 3834
rect 11236 3782 11238 3834
rect 11238 3782 11290 3834
rect 11290 3782 11292 3834
rect 10916 3780 10972 3782
rect 10996 3780 11052 3782
rect 11076 3780 11132 3782
rect 11156 3780 11212 3782
rect 11236 3780 11292 3782
rect 11656 3290 11712 3292
rect 11736 3290 11792 3292
rect 11816 3290 11872 3292
rect 11896 3290 11952 3292
rect 11976 3290 12032 3292
rect 11656 3238 11658 3290
rect 11658 3238 11710 3290
rect 11710 3238 11712 3290
rect 11736 3238 11774 3290
rect 11774 3238 11786 3290
rect 11786 3238 11792 3290
rect 11816 3238 11838 3290
rect 11838 3238 11850 3290
rect 11850 3238 11872 3290
rect 11896 3238 11902 3290
rect 11902 3238 11914 3290
rect 11914 3238 11952 3290
rect 11976 3238 11978 3290
rect 11978 3238 12030 3290
rect 12030 3238 12032 3290
rect 11656 3236 11712 3238
rect 11736 3236 11792 3238
rect 11816 3236 11872 3238
rect 11896 3236 11952 3238
rect 11976 3236 12032 3238
rect 14916 10362 14972 10364
rect 14996 10362 15052 10364
rect 15076 10362 15132 10364
rect 15156 10362 15212 10364
rect 15236 10362 15292 10364
rect 14916 10310 14918 10362
rect 14918 10310 14970 10362
rect 14970 10310 14972 10362
rect 14996 10310 15034 10362
rect 15034 10310 15046 10362
rect 15046 10310 15052 10362
rect 15076 10310 15098 10362
rect 15098 10310 15110 10362
rect 15110 10310 15132 10362
rect 15156 10310 15162 10362
rect 15162 10310 15174 10362
rect 15174 10310 15212 10362
rect 15236 10310 15238 10362
rect 15238 10310 15290 10362
rect 15290 10310 15292 10362
rect 14916 10308 14972 10310
rect 14996 10308 15052 10310
rect 15076 10308 15132 10310
rect 15156 10308 15212 10310
rect 15236 10308 15292 10310
rect 15656 15258 15712 15260
rect 15736 15258 15792 15260
rect 15816 15258 15872 15260
rect 15896 15258 15952 15260
rect 15976 15258 16032 15260
rect 15656 15206 15658 15258
rect 15658 15206 15710 15258
rect 15710 15206 15712 15258
rect 15736 15206 15774 15258
rect 15774 15206 15786 15258
rect 15786 15206 15792 15258
rect 15816 15206 15838 15258
rect 15838 15206 15850 15258
rect 15850 15206 15872 15258
rect 15896 15206 15902 15258
rect 15902 15206 15914 15258
rect 15914 15206 15952 15258
rect 15976 15206 15978 15258
rect 15978 15206 16030 15258
rect 16030 15206 16032 15258
rect 15656 15204 15712 15206
rect 15736 15204 15792 15206
rect 15816 15204 15872 15206
rect 15896 15204 15952 15206
rect 15976 15204 16032 15206
rect 15750 14456 15806 14512
rect 15656 14170 15712 14172
rect 15736 14170 15792 14172
rect 15816 14170 15872 14172
rect 15896 14170 15952 14172
rect 15976 14170 16032 14172
rect 15656 14118 15658 14170
rect 15658 14118 15710 14170
rect 15710 14118 15712 14170
rect 15736 14118 15774 14170
rect 15774 14118 15786 14170
rect 15786 14118 15792 14170
rect 15816 14118 15838 14170
rect 15838 14118 15850 14170
rect 15850 14118 15872 14170
rect 15896 14118 15902 14170
rect 15902 14118 15914 14170
rect 15914 14118 15952 14170
rect 15976 14118 15978 14170
rect 15978 14118 16030 14170
rect 16030 14118 16032 14170
rect 15656 14116 15712 14118
rect 15736 14116 15792 14118
rect 15816 14116 15872 14118
rect 15896 14116 15952 14118
rect 15976 14116 16032 14118
rect 15656 13082 15712 13084
rect 15736 13082 15792 13084
rect 15816 13082 15872 13084
rect 15896 13082 15952 13084
rect 15976 13082 16032 13084
rect 15656 13030 15658 13082
rect 15658 13030 15710 13082
rect 15710 13030 15712 13082
rect 15736 13030 15774 13082
rect 15774 13030 15786 13082
rect 15786 13030 15792 13082
rect 15816 13030 15838 13082
rect 15838 13030 15850 13082
rect 15850 13030 15872 13082
rect 15896 13030 15902 13082
rect 15902 13030 15914 13082
rect 15914 13030 15952 13082
rect 15976 13030 15978 13082
rect 15978 13030 16030 13082
rect 16030 13030 16032 13082
rect 15656 13028 15712 13030
rect 15736 13028 15792 13030
rect 15816 13028 15872 13030
rect 15896 13028 15952 13030
rect 15976 13028 16032 13030
rect 15656 11994 15712 11996
rect 15736 11994 15792 11996
rect 15816 11994 15872 11996
rect 15896 11994 15952 11996
rect 15976 11994 16032 11996
rect 15656 11942 15658 11994
rect 15658 11942 15710 11994
rect 15710 11942 15712 11994
rect 15736 11942 15774 11994
rect 15774 11942 15786 11994
rect 15786 11942 15792 11994
rect 15816 11942 15838 11994
rect 15838 11942 15850 11994
rect 15850 11942 15872 11994
rect 15896 11942 15902 11994
rect 15902 11942 15914 11994
rect 15914 11942 15952 11994
rect 15976 11942 15978 11994
rect 15978 11942 16030 11994
rect 16030 11942 16032 11994
rect 15656 11940 15712 11942
rect 15736 11940 15792 11942
rect 15816 11940 15872 11942
rect 15896 11940 15952 11942
rect 15976 11940 16032 11942
rect 15656 10906 15712 10908
rect 15736 10906 15792 10908
rect 15816 10906 15872 10908
rect 15896 10906 15952 10908
rect 15976 10906 16032 10908
rect 15656 10854 15658 10906
rect 15658 10854 15710 10906
rect 15710 10854 15712 10906
rect 15736 10854 15774 10906
rect 15774 10854 15786 10906
rect 15786 10854 15792 10906
rect 15816 10854 15838 10906
rect 15838 10854 15850 10906
rect 15850 10854 15872 10906
rect 15896 10854 15902 10906
rect 15902 10854 15914 10906
rect 15914 10854 15952 10906
rect 15976 10854 15978 10906
rect 15978 10854 16030 10906
rect 16030 10854 16032 10906
rect 15656 10852 15712 10854
rect 15736 10852 15792 10854
rect 15816 10852 15872 10854
rect 15896 10852 15952 10854
rect 15976 10852 16032 10854
rect 17682 24928 17738 24984
rect 16578 22480 16634 22536
rect 16578 15952 16634 16008
rect 15656 9818 15712 9820
rect 15736 9818 15792 9820
rect 15816 9818 15872 9820
rect 15896 9818 15952 9820
rect 15976 9818 16032 9820
rect 15656 9766 15658 9818
rect 15658 9766 15710 9818
rect 15710 9766 15712 9818
rect 15736 9766 15774 9818
rect 15774 9766 15786 9818
rect 15786 9766 15792 9818
rect 15816 9766 15838 9818
rect 15838 9766 15850 9818
rect 15850 9766 15872 9818
rect 15896 9766 15902 9818
rect 15902 9766 15914 9818
rect 15914 9766 15952 9818
rect 15976 9766 15978 9818
rect 15978 9766 16030 9818
rect 16030 9766 16032 9818
rect 15656 9764 15712 9766
rect 15736 9764 15792 9766
rect 15816 9764 15872 9766
rect 15896 9764 15952 9766
rect 15976 9764 16032 9766
rect 14916 9274 14972 9276
rect 14996 9274 15052 9276
rect 15076 9274 15132 9276
rect 15156 9274 15212 9276
rect 15236 9274 15292 9276
rect 14916 9222 14918 9274
rect 14918 9222 14970 9274
rect 14970 9222 14972 9274
rect 14996 9222 15034 9274
rect 15034 9222 15046 9274
rect 15046 9222 15052 9274
rect 15076 9222 15098 9274
rect 15098 9222 15110 9274
rect 15110 9222 15132 9274
rect 15156 9222 15162 9274
rect 15162 9222 15174 9274
rect 15174 9222 15212 9274
rect 15236 9222 15238 9274
rect 15238 9222 15290 9274
rect 15290 9222 15292 9274
rect 14916 9220 14972 9222
rect 14996 9220 15052 9222
rect 15076 9220 15132 9222
rect 15156 9220 15212 9222
rect 15236 9220 15292 9222
rect 14916 8186 14972 8188
rect 14996 8186 15052 8188
rect 15076 8186 15132 8188
rect 15156 8186 15212 8188
rect 15236 8186 15292 8188
rect 14916 8134 14918 8186
rect 14918 8134 14970 8186
rect 14970 8134 14972 8186
rect 14996 8134 15034 8186
rect 15034 8134 15046 8186
rect 15046 8134 15052 8186
rect 15076 8134 15098 8186
rect 15098 8134 15110 8186
rect 15110 8134 15132 8186
rect 15156 8134 15162 8186
rect 15162 8134 15174 8186
rect 15174 8134 15212 8186
rect 15236 8134 15238 8186
rect 15238 8134 15290 8186
rect 15290 8134 15292 8186
rect 14916 8132 14972 8134
rect 14996 8132 15052 8134
rect 15076 8132 15132 8134
rect 15156 8132 15212 8134
rect 15236 8132 15292 8134
rect 15656 8730 15712 8732
rect 15736 8730 15792 8732
rect 15816 8730 15872 8732
rect 15896 8730 15952 8732
rect 15976 8730 16032 8732
rect 15656 8678 15658 8730
rect 15658 8678 15710 8730
rect 15710 8678 15712 8730
rect 15736 8678 15774 8730
rect 15774 8678 15786 8730
rect 15786 8678 15792 8730
rect 15816 8678 15838 8730
rect 15838 8678 15850 8730
rect 15850 8678 15872 8730
rect 15896 8678 15902 8730
rect 15902 8678 15914 8730
rect 15914 8678 15952 8730
rect 15976 8678 15978 8730
rect 15978 8678 16030 8730
rect 16030 8678 16032 8730
rect 15656 8676 15712 8678
rect 15736 8676 15792 8678
rect 15816 8676 15872 8678
rect 15896 8676 15952 8678
rect 15976 8676 16032 8678
rect 15382 7792 15438 7848
rect 14916 7098 14972 7100
rect 14996 7098 15052 7100
rect 15076 7098 15132 7100
rect 15156 7098 15212 7100
rect 15236 7098 15292 7100
rect 14916 7046 14918 7098
rect 14918 7046 14970 7098
rect 14970 7046 14972 7098
rect 14996 7046 15034 7098
rect 15034 7046 15046 7098
rect 15046 7046 15052 7098
rect 15076 7046 15098 7098
rect 15098 7046 15110 7098
rect 15110 7046 15132 7098
rect 15156 7046 15162 7098
rect 15162 7046 15174 7098
rect 15174 7046 15212 7098
rect 15236 7046 15238 7098
rect 15238 7046 15290 7098
rect 15290 7046 15292 7098
rect 14916 7044 14972 7046
rect 14996 7044 15052 7046
rect 15076 7044 15132 7046
rect 15156 7044 15212 7046
rect 15236 7044 15292 7046
rect 15656 7642 15712 7644
rect 15736 7642 15792 7644
rect 15816 7642 15872 7644
rect 15896 7642 15952 7644
rect 15976 7642 16032 7644
rect 15656 7590 15658 7642
rect 15658 7590 15710 7642
rect 15710 7590 15712 7642
rect 15736 7590 15774 7642
rect 15774 7590 15786 7642
rect 15786 7590 15792 7642
rect 15816 7590 15838 7642
rect 15838 7590 15850 7642
rect 15850 7590 15872 7642
rect 15896 7590 15902 7642
rect 15902 7590 15914 7642
rect 15914 7590 15952 7642
rect 15976 7590 15978 7642
rect 15978 7590 16030 7642
rect 16030 7590 16032 7642
rect 15656 7588 15712 7590
rect 15736 7588 15792 7590
rect 15816 7588 15872 7590
rect 15896 7588 15952 7590
rect 15976 7588 16032 7590
rect 15656 6554 15712 6556
rect 15736 6554 15792 6556
rect 15816 6554 15872 6556
rect 15896 6554 15952 6556
rect 15976 6554 16032 6556
rect 15656 6502 15658 6554
rect 15658 6502 15710 6554
rect 15710 6502 15712 6554
rect 15736 6502 15774 6554
rect 15774 6502 15786 6554
rect 15786 6502 15792 6554
rect 15816 6502 15838 6554
rect 15838 6502 15850 6554
rect 15850 6502 15872 6554
rect 15896 6502 15902 6554
rect 15902 6502 15914 6554
rect 15914 6502 15952 6554
rect 15976 6502 15978 6554
rect 15978 6502 16030 6554
rect 16030 6502 16032 6554
rect 15656 6500 15712 6502
rect 15736 6500 15792 6502
rect 15816 6500 15872 6502
rect 15896 6500 15952 6502
rect 15976 6500 16032 6502
rect 14916 6010 14972 6012
rect 14996 6010 15052 6012
rect 15076 6010 15132 6012
rect 15156 6010 15212 6012
rect 15236 6010 15292 6012
rect 14916 5958 14918 6010
rect 14918 5958 14970 6010
rect 14970 5958 14972 6010
rect 14996 5958 15034 6010
rect 15034 5958 15046 6010
rect 15046 5958 15052 6010
rect 15076 5958 15098 6010
rect 15098 5958 15110 6010
rect 15110 5958 15132 6010
rect 15156 5958 15162 6010
rect 15162 5958 15174 6010
rect 15174 5958 15212 6010
rect 15236 5958 15238 6010
rect 15238 5958 15290 6010
rect 15290 5958 15292 6010
rect 14916 5956 14972 5958
rect 14996 5956 15052 5958
rect 15076 5956 15132 5958
rect 15156 5956 15212 5958
rect 15236 5956 15292 5958
rect 15656 5466 15712 5468
rect 15736 5466 15792 5468
rect 15816 5466 15872 5468
rect 15896 5466 15952 5468
rect 15976 5466 16032 5468
rect 15656 5414 15658 5466
rect 15658 5414 15710 5466
rect 15710 5414 15712 5466
rect 15736 5414 15774 5466
rect 15774 5414 15786 5466
rect 15786 5414 15792 5466
rect 15816 5414 15838 5466
rect 15838 5414 15850 5466
rect 15850 5414 15872 5466
rect 15896 5414 15902 5466
rect 15902 5414 15914 5466
rect 15914 5414 15952 5466
rect 15976 5414 15978 5466
rect 15978 5414 16030 5466
rect 16030 5414 16032 5466
rect 15656 5412 15712 5414
rect 15736 5412 15792 5414
rect 15816 5412 15872 5414
rect 15896 5412 15952 5414
rect 15976 5412 16032 5414
rect 6916 2746 6972 2748
rect 6996 2746 7052 2748
rect 7076 2746 7132 2748
rect 7156 2746 7212 2748
rect 7236 2746 7292 2748
rect 6916 2694 6918 2746
rect 6918 2694 6970 2746
rect 6970 2694 6972 2746
rect 6996 2694 7034 2746
rect 7034 2694 7046 2746
rect 7046 2694 7052 2746
rect 7076 2694 7098 2746
rect 7098 2694 7110 2746
rect 7110 2694 7132 2746
rect 7156 2694 7162 2746
rect 7162 2694 7174 2746
rect 7174 2694 7212 2746
rect 7236 2694 7238 2746
rect 7238 2694 7290 2746
rect 7290 2694 7292 2746
rect 6916 2692 6972 2694
rect 6996 2692 7052 2694
rect 7076 2692 7132 2694
rect 7156 2692 7212 2694
rect 7236 2692 7292 2694
rect 14916 4922 14972 4924
rect 14996 4922 15052 4924
rect 15076 4922 15132 4924
rect 15156 4922 15212 4924
rect 15236 4922 15292 4924
rect 14916 4870 14918 4922
rect 14918 4870 14970 4922
rect 14970 4870 14972 4922
rect 14996 4870 15034 4922
rect 15034 4870 15046 4922
rect 15046 4870 15052 4922
rect 15076 4870 15098 4922
rect 15098 4870 15110 4922
rect 15110 4870 15132 4922
rect 15156 4870 15162 4922
rect 15162 4870 15174 4922
rect 15174 4870 15212 4922
rect 15236 4870 15238 4922
rect 15238 4870 15290 4922
rect 15290 4870 15292 4922
rect 14916 4868 14972 4870
rect 14996 4868 15052 4870
rect 15076 4868 15132 4870
rect 15156 4868 15212 4870
rect 15236 4868 15292 4870
rect 15656 4378 15712 4380
rect 15736 4378 15792 4380
rect 15816 4378 15872 4380
rect 15896 4378 15952 4380
rect 15976 4378 16032 4380
rect 15656 4326 15658 4378
rect 15658 4326 15710 4378
rect 15710 4326 15712 4378
rect 15736 4326 15774 4378
rect 15774 4326 15786 4378
rect 15786 4326 15792 4378
rect 15816 4326 15838 4378
rect 15838 4326 15850 4378
rect 15850 4326 15872 4378
rect 15896 4326 15902 4378
rect 15902 4326 15914 4378
rect 15914 4326 15952 4378
rect 15976 4326 15978 4378
rect 15978 4326 16030 4378
rect 16030 4326 16032 4378
rect 15656 4324 15712 4326
rect 15736 4324 15792 4326
rect 15816 4324 15872 4326
rect 15896 4324 15952 4326
rect 15976 4324 16032 4326
rect 17590 18128 17646 18184
rect 17774 16224 17830 16280
rect 19656 27226 19712 27228
rect 19736 27226 19792 27228
rect 19816 27226 19872 27228
rect 19896 27226 19952 27228
rect 19976 27226 20032 27228
rect 19656 27174 19658 27226
rect 19658 27174 19710 27226
rect 19710 27174 19712 27226
rect 19736 27174 19774 27226
rect 19774 27174 19786 27226
rect 19786 27174 19792 27226
rect 19816 27174 19838 27226
rect 19838 27174 19850 27226
rect 19850 27174 19872 27226
rect 19896 27174 19902 27226
rect 19902 27174 19914 27226
rect 19914 27174 19952 27226
rect 19976 27174 19978 27226
rect 19978 27174 20030 27226
rect 20030 27174 20032 27226
rect 19656 27172 19712 27174
rect 19736 27172 19792 27174
rect 19816 27172 19872 27174
rect 19896 27172 19952 27174
rect 19976 27172 20032 27174
rect 18916 26682 18972 26684
rect 18996 26682 19052 26684
rect 19076 26682 19132 26684
rect 19156 26682 19212 26684
rect 19236 26682 19292 26684
rect 18916 26630 18918 26682
rect 18918 26630 18970 26682
rect 18970 26630 18972 26682
rect 18996 26630 19034 26682
rect 19034 26630 19046 26682
rect 19046 26630 19052 26682
rect 19076 26630 19098 26682
rect 19098 26630 19110 26682
rect 19110 26630 19132 26682
rect 19156 26630 19162 26682
rect 19162 26630 19174 26682
rect 19174 26630 19212 26682
rect 19236 26630 19238 26682
rect 19238 26630 19290 26682
rect 19290 26630 19292 26682
rect 18916 26628 18972 26630
rect 18996 26628 19052 26630
rect 19076 26628 19132 26630
rect 19156 26628 19212 26630
rect 19236 26628 19292 26630
rect 18916 25594 18972 25596
rect 18996 25594 19052 25596
rect 19076 25594 19132 25596
rect 19156 25594 19212 25596
rect 19236 25594 19292 25596
rect 18916 25542 18918 25594
rect 18918 25542 18970 25594
rect 18970 25542 18972 25594
rect 18996 25542 19034 25594
rect 19034 25542 19046 25594
rect 19046 25542 19052 25594
rect 19076 25542 19098 25594
rect 19098 25542 19110 25594
rect 19110 25542 19132 25594
rect 19156 25542 19162 25594
rect 19162 25542 19174 25594
rect 19174 25542 19212 25594
rect 19236 25542 19238 25594
rect 19238 25542 19290 25594
rect 19290 25542 19292 25594
rect 18916 25540 18972 25542
rect 18996 25540 19052 25542
rect 19076 25540 19132 25542
rect 19156 25540 19212 25542
rect 19236 25540 19292 25542
rect 19656 26138 19712 26140
rect 19736 26138 19792 26140
rect 19816 26138 19872 26140
rect 19896 26138 19952 26140
rect 19976 26138 20032 26140
rect 19656 26086 19658 26138
rect 19658 26086 19710 26138
rect 19710 26086 19712 26138
rect 19736 26086 19774 26138
rect 19774 26086 19786 26138
rect 19786 26086 19792 26138
rect 19816 26086 19838 26138
rect 19838 26086 19850 26138
rect 19850 26086 19872 26138
rect 19896 26086 19902 26138
rect 19902 26086 19914 26138
rect 19914 26086 19952 26138
rect 19976 26086 19978 26138
rect 19978 26086 20030 26138
rect 20030 26086 20032 26138
rect 19656 26084 19712 26086
rect 19736 26084 19792 26086
rect 19816 26084 19872 26086
rect 19896 26084 19952 26086
rect 19976 26084 20032 26086
rect 19656 25050 19712 25052
rect 19736 25050 19792 25052
rect 19816 25050 19872 25052
rect 19896 25050 19952 25052
rect 19976 25050 20032 25052
rect 19656 24998 19658 25050
rect 19658 24998 19710 25050
rect 19710 24998 19712 25050
rect 19736 24998 19774 25050
rect 19774 24998 19786 25050
rect 19786 24998 19792 25050
rect 19816 24998 19838 25050
rect 19838 24998 19850 25050
rect 19850 24998 19872 25050
rect 19896 24998 19902 25050
rect 19902 24998 19914 25050
rect 19914 24998 19952 25050
rect 19976 24998 19978 25050
rect 19978 24998 20030 25050
rect 20030 24998 20032 25050
rect 19656 24996 19712 24998
rect 19736 24996 19792 24998
rect 19816 24996 19872 24998
rect 19896 24996 19952 24998
rect 19976 24996 20032 24998
rect 18916 24506 18972 24508
rect 18996 24506 19052 24508
rect 19076 24506 19132 24508
rect 19156 24506 19212 24508
rect 19236 24506 19292 24508
rect 18916 24454 18918 24506
rect 18918 24454 18970 24506
rect 18970 24454 18972 24506
rect 18996 24454 19034 24506
rect 19034 24454 19046 24506
rect 19046 24454 19052 24506
rect 19076 24454 19098 24506
rect 19098 24454 19110 24506
rect 19110 24454 19132 24506
rect 19156 24454 19162 24506
rect 19162 24454 19174 24506
rect 19174 24454 19212 24506
rect 19236 24454 19238 24506
rect 19238 24454 19290 24506
rect 19290 24454 19292 24506
rect 18916 24452 18972 24454
rect 18996 24452 19052 24454
rect 19076 24452 19132 24454
rect 19156 24452 19212 24454
rect 19236 24452 19292 24454
rect 18916 23418 18972 23420
rect 18996 23418 19052 23420
rect 19076 23418 19132 23420
rect 19156 23418 19212 23420
rect 19236 23418 19292 23420
rect 18916 23366 18918 23418
rect 18918 23366 18970 23418
rect 18970 23366 18972 23418
rect 18996 23366 19034 23418
rect 19034 23366 19046 23418
rect 19046 23366 19052 23418
rect 19076 23366 19098 23418
rect 19098 23366 19110 23418
rect 19110 23366 19132 23418
rect 19156 23366 19162 23418
rect 19162 23366 19174 23418
rect 19174 23366 19212 23418
rect 19236 23366 19238 23418
rect 19238 23366 19290 23418
rect 19290 23366 19292 23418
rect 18916 23364 18972 23366
rect 18996 23364 19052 23366
rect 19076 23364 19132 23366
rect 19156 23364 19212 23366
rect 19236 23364 19292 23366
rect 19656 23962 19712 23964
rect 19736 23962 19792 23964
rect 19816 23962 19872 23964
rect 19896 23962 19952 23964
rect 19976 23962 20032 23964
rect 19656 23910 19658 23962
rect 19658 23910 19710 23962
rect 19710 23910 19712 23962
rect 19736 23910 19774 23962
rect 19774 23910 19786 23962
rect 19786 23910 19792 23962
rect 19816 23910 19838 23962
rect 19838 23910 19850 23962
rect 19850 23910 19872 23962
rect 19896 23910 19902 23962
rect 19902 23910 19914 23962
rect 19914 23910 19952 23962
rect 19976 23910 19978 23962
rect 19978 23910 20030 23962
rect 20030 23910 20032 23962
rect 19656 23908 19712 23910
rect 19736 23908 19792 23910
rect 19816 23908 19872 23910
rect 19896 23908 19952 23910
rect 19976 23908 20032 23910
rect 18916 22330 18972 22332
rect 18996 22330 19052 22332
rect 19076 22330 19132 22332
rect 19156 22330 19212 22332
rect 19236 22330 19292 22332
rect 18916 22278 18918 22330
rect 18918 22278 18970 22330
rect 18970 22278 18972 22330
rect 18996 22278 19034 22330
rect 19034 22278 19046 22330
rect 19046 22278 19052 22330
rect 19076 22278 19098 22330
rect 19098 22278 19110 22330
rect 19110 22278 19132 22330
rect 19156 22278 19162 22330
rect 19162 22278 19174 22330
rect 19174 22278 19212 22330
rect 19236 22278 19238 22330
rect 19238 22278 19290 22330
rect 19290 22278 19292 22330
rect 18916 22276 18972 22278
rect 18996 22276 19052 22278
rect 19076 22276 19132 22278
rect 19156 22276 19212 22278
rect 19236 22276 19292 22278
rect 19890 23060 19892 23080
rect 19892 23060 19944 23080
rect 19944 23060 19946 23080
rect 19890 23024 19946 23060
rect 19656 22874 19712 22876
rect 19736 22874 19792 22876
rect 19816 22874 19872 22876
rect 19896 22874 19952 22876
rect 19976 22874 20032 22876
rect 19656 22822 19658 22874
rect 19658 22822 19710 22874
rect 19710 22822 19712 22874
rect 19736 22822 19774 22874
rect 19774 22822 19786 22874
rect 19786 22822 19792 22874
rect 19816 22822 19838 22874
rect 19838 22822 19850 22874
rect 19850 22822 19872 22874
rect 19896 22822 19902 22874
rect 19902 22822 19914 22874
rect 19914 22822 19952 22874
rect 19976 22822 19978 22874
rect 19978 22822 20030 22874
rect 20030 22822 20032 22874
rect 19656 22820 19712 22822
rect 19736 22820 19792 22822
rect 19816 22820 19872 22822
rect 19896 22820 19952 22822
rect 19976 22820 20032 22822
rect 19890 22616 19946 22672
rect 19890 22072 19946 22128
rect 18916 21242 18972 21244
rect 18996 21242 19052 21244
rect 19076 21242 19132 21244
rect 19156 21242 19212 21244
rect 19236 21242 19292 21244
rect 18916 21190 18918 21242
rect 18918 21190 18970 21242
rect 18970 21190 18972 21242
rect 18996 21190 19034 21242
rect 19034 21190 19046 21242
rect 19046 21190 19052 21242
rect 19076 21190 19098 21242
rect 19098 21190 19110 21242
rect 19110 21190 19132 21242
rect 19156 21190 19162 21242
rect 19162 21190 19174 21242
rect 19174 21190 19212 21242
rect 19236 21190 19238 21242
rect 19238 21190 19290 21242
rect 19290 21190 19292 21242
rect 18916 21188 18972 21190
rect 18996 21188 19052 21190
rect 19076 21188 19132 21190
rect 19156 21188 19212 21190
rect 19236 21188 19292 21190
rect 18326 20340 18328 20360
rect 18328 20340 18380 20360
rect 18380 20340 18382 20360
rect 18326 20304 18382 20340
rect 19656 21786 19712 21788
rect 19736 21786 19792 21788
rect 19816 21786 19872 21788
rect 19896 21786 19952 21788
rect 19976 21786 20032 21788
rect 19656 21734 19658 21786
rect 19658 21734 19710 21786
rect 19710 21734 19712 21786
rect 19736 21734 19774 21786
rect 19774 21734 19786 21786
rect 19786 21734 19792 21786
rect 19816 21734 19838 21786
rect 19838 21734 19850 21786
rect 19850 21734 19872 21786
rect 19896 21734 19902 21786
rect 19902 21734 19914 21786
rect 19914 21734 19952 21786
rect 19976 21734 19978 21786
rect 19978 21734 20030 21786
rect 20030 21734 20032 21786
rect 19656 21732 19712 21734
rect 19736 21732 19792 21734
rect 19816 21732 19872 21734
rect 19896 21732 19952 21734
rect 19976 21732 20032 21734
rect 19614 20848 19670 20904
rect 19656 20698 19712 20700
rect 19736 20698 19792 20700
rect 19816 20698 19872 20700
rect 19896 20698 19952 20700
rect 19976 20698 20032 20700
rect 19656 20646 19658 20698
rect 19658 20646 19710 20698
rect 19710 20646 19712 20698
rect 19736 20646 19774 20698
rect 19774 20646 19786 20698
rect 19786 20646 19792 20698
rect 19816 20646 19838 20698
rect 19838 20646 19850 20698
rect 19850 20646 19872 20698
rect 19896 20646 19902 20698
rect 19902 20646 19914 20698
rect 19914 20646 19952 20698
rect 19976 20646 19978 20698
rect 19978 20646 20030 20698
rect 20030 20646 20032 20698
rect 19656 20644 19712 20646
rect 19736 20644 19792 20646
rect 19816 20644 19872 20646
rect 19896 20644 19952 20646
rect 19976 20644 20032 20646
rect 17314 10668 17370 10704
rect 17314 10648 17316 10668
rect 17316 10648 17368 10668
rect 17368 10648 17370 10668
rect 14916 3834 14972 3836
rect 14996 3834 15052 3836
rect 15076 3834 15132 3836
rect 15156 3834 15212 3836
rect 15236 3834 15292 3836
rect 14916 3782 14918 3834
rect 14918 3782 14970 3834
rect 14970 3782 14972 3834
rect 14996 3782 15034 3834
rect 15034 3782 15046 3834
rect 15046 3782 15052 3834
rect 15076 3782 15098 3834
rect 15098 3782 15110 3834
rect 15110 3782 15132 3834
rect 15156 3782 15162 3834
rect 15162 3782 15174 3834
rect 15174 3782 15212 3834
rect 15236 3782 15238 3834
rect 15238 3782 15290 3834
rect 15290 3782 15292 3834
rect 14916 3780 14972 3782
rect 14996 3780 15052 3782
rect 15076 3780 15132 3782
rect 15156 3780 15212 3782
rect 15236 3780 15292 3782
rect 15656 3290 15712 3292
rect 15736 3290 15792 3292
rect 15816 3290 15872 3292
rect 15896 3290 15952 3292
rect 15976 3290 16032 3292
rect 15656 3238 15658 3290
rect 15658 3238 15710 3290
rect 15710 3238 15712 3290
rect 15736 3238 15774 3290
rect 15774 3238 15786 3290
rect 15786 3238 15792 3290
rect 15816 3238 15838 3290
rect 15838 3238 15850 3290
rect 15850 3238 15872 3290
rect 15896 3238 15902 3290
rect 15902 3238 15914 3290
rect 15914 3238 15952 3290
rect 15976 3238 15978 3290
rect 15978 3238 16030 3290
rect 16030 3238 16032 3290
rect 15656 3236 15712 3238
rect 15736 3236 15792 3238
rect 15816 3236 15872 3238
rect 15896 3236 15952 3238
rect 15976 3236 16032 3238
rect 17498 10260 17554 10296
rect 17498 10240 17500 10260
rect 17500 10240 17552 10260
rect 17552 10240 17554 10260
rect 17590 9968 17646 10024
rect 18234 15408 18290 15464
rect 18050 6704 18106 6760
rect 18602 17040 18658 17096
rect 18916 20154 18972 20156
rect 18996 20154 19052 20156
rect 19076 20154 19132 20156
rect 19156 20154 19212 20156
rect 19236 20154 19292 20156
rect 18916 20102 18918 20154
rect 18918 20102 18970 20154
rect 18970 20102 18972 20154
rect 18996 20102 19034 20154
rect 19034 20102 19046 20154
rect 19046 20102 19052 20154
rect 19076 20102 19098 20154
rect 19098 20102 19110 20154
rect 19110 20102 19132 20154
rect 19156 20102 19162 20154
rect 19162 20102 19174 20154
rect 19174 20102 19212 20154
rect 19236 20102 19238 20154
rect 19238 20102 19290 20154
rect 19290 20102 19292 20154
rect 18916 20100 18972 20102
rect 18996 20100 19052 20102
rect 19076 20100 19132 20102
rect 19156 20100 19212 20102
rect 19236 20100 19292 20102
rect 18916 19066 18972 19068
rect 18996 19066 19052 19068
rect 19076 19066 19132 19068
rect 19156 19066 19212 19068
rect 19236 19066 19292 19068
rect 18916 19014 18918 19066
rect 18918 19014 18970 19066
rect 18970 19014 18972 19066
rect 18996 19014 19034 19066
rect 19034 19014 19046 19066
rect 19046 19014 19052 19066
rect 19076 19014 19098 19066
rect 19098 19014 19110 19066
rect 19110 19014 19132 19066
rect 19156 19014 19162 19066
rect 19162 19014 19174 19066
rect 19174 19014 19212 19066
rect 19236 19014 19238 19066
rect 19238 19014 19290 19066
rect 19290 19014 19292 19066
rect 18916 19012 18972 19014
rect 18996 19012 19052 19014
rect 19076 19012 19132 19014
rect 19156 19012 19212 19014
rect 19236 19012 19292 19014
rect 19656 19610 19712 19612
rect 19736 19610 19792 19612
rect 19816 19610 19872 19612
rect 19896 19610 19952 19612
rect 19976 19610 20032 19612
rect 19656 19558 19658 19610
rect 19658 19558 19710 19610
rect 19710 19558 19712 19610
rect 19736 19558 19774 19610
rect 19774 19558 19786 19610
rect 19786 19558 19792 19610
rect 19816 19558 19838 19610
rect 19838 19558 19850 19610
rect 19850 19558 19872 19610
rect 19896 19558 19902 19610
rect 19902 19558 19914 19610
rect 19914 19558 19952 19610
rect 19976 19558 19978 19610
rect 19978 19558 20030 19610
rect 20030 19558 20032 19610
rect 19656 19556 19712 19558
rect 19736 19556 19792 19558
rect 19816 19556 19872 19558
rect 19896 19556 19952 19558
rect 19976 19556 20032 19558
rect 20534 21936 20590 21992
rect 19656 18522 19712 18524
rect 19736 18522 19792 18524
rect 19816 18522 19872 18524
rect 19896 18522 19952 18524
rect 19976 18522 20032 18524
rect 19656 18470 19658 18522
rect 19658 18470 19710 18522
rect 19710 18470 19712 18522
rect 19736 18470 19774 18522
rect 19774 18470 19786 18522
rect 19786 18470 19792 18522
rect 19816 18470 19838 18522
rect 19838 18470 19850 18522
rect 19850 18470 19872 18522
rect 19896 18470 19902 18522
rect 19902 18470 19914 18522
rect 19914 18470 19952 18522
rect 19976 18470 19978 18522
rect 19978 18470 20030 18522
rect 20030 18470 20032 18522
rect 19656 18468 19712 18470
rect 19736 18468 19792 18470
rect 19816 18468 19872 18470
rect 19896 18468 19952 18470
rect 19976 18468 20032 18470
rect 18916 17978 18972 17980
rect 18996 17978 19052 17980
rect 19076 17978 19132 17980
rect 19156 17978 19212 17980
rect 19236 17978 19292 17980
rect 18916 17926 18918 17978
rect 18918 17926 18970 17978
rect 18970 17926 18972 17978
rect 18996 17926 19034 17978
rect 19034 17926 19046 17978
rect 19046 17926 19052 17978
rect 19076 17926 19098 17978
rect 19098 17926 19110 17978
rect 19110 17926 19132 17978
rect 19156 17926 19162 17978
rect 19162 17926 19174 17978
rect 19174 17926 19212 17978
rect 19236 17926 19238 17978
rect 19238 17926 19290 17978
rect 19290 17926 19292 17978
rect 18916 17924 18972 17926
rect 18996 17924 19052 17926
rect 19076 17924 19132 17926
rect 19156 17924 19212 17926
rect 19236 17924 19292 17926
rect 19656 17434 19712 17436
rect 19736 17434 19792 17436
rect 19816 17434 19872 17436
rect 19896 17434 19952 17436
rect 19976 17434 20032 17436
rect 19656 17382 19658 17434
rect 19658 17382 19710 17434
rect 19710 17382 19712 17434
rect 19736 17382 19774 17434
rect 19774 17382 19786 17434
rect 19786 17382 19792 17434
rect 19816 17382 19838 17434
rect 19838 17382 19850 17434
rect 19850 17382 19872 17434
rect 19896 17382 19902 17434
rect 19902 17382 19914 17434
rect 19914 17382 19952 17434
rect 19976 17382 19978 17434
rect 19978 17382 20030 17434
rect 20030 17382 20032 17434
rect 19656 17380 19712 17382
rect 19736 17380 19792 17382
rect 19816 17380 19872 17382
rect 19896 17380 19952 17382
rect 19976 17380 20032 17382
rect 18916 16890 18972 16892
rect 18996 16890 19052 16892
rect 19076 16890 19132 16892
rect 19156 16890 19212 16892
rect 19236 16890 19292 16892
rect 18916 16838 18918 16890
rect 18918 16838 18970 16890
rect 18970 16838 18972 16890
rect 18996 16838 19034 16890
rect 19034 16838 19046 16890
rect 19046 16838 19052 16890
rect 19076 16838 19098 16890
rect 19098 16838 19110 16890
rect 19110 16838 19132 16890
rect 19156 16838 19162 16890
rect 19162 16838 19174 16890
rect 19174 16838 19212 16890
rect 19236 16838 19238 16890
rect 19238 16838 19290 16890
rect 19290 16838 19292 16890
rect 18916 16836 18972 16838
rect 18996 16836 19052 16838
rect 19076 16836 19132 16838
rect 19156 16836 19212 16838
rect 19236 16836 19292 16838
rect 18970 16496 19026 16552
rect 18786 16224 18842 16280
rect 19338 16244 19394 16280
rect 19338 16224 19340 16244
rect 19340 16224 19392 16244
rect 19392 16224 19394 16244
rect 18916 15802 18972 15804
rect 18996 15802 19052 15804
rect 19076 15802 19132 15804
rect 19156 15802 19212 15804
rect 19236 15802 19292 15804
rect 18916 15750 18918 15802
rect 18918 15750 18970 15802
rect 18970 15750 18972 15802
rect 18996 15750 19034 15802
rect 19034 15750 19046 15802
rect 19046 15750 19052 15802
rect 19076 15750 19098 15802
rect 19098 15750 19110 15802
rect 19110 15750 19132 15802
rect 19156 15750 19162 15802
rect 19162 15750 19174 15802
rect 19174 15750 19212 15802
rect 19236 15750 19238 15802
rect 19238 15750 19290 15802
rect 19290 15750 19292 15802
rect 18916 15748 18972 15750
rect 18996 15748 19052 15750
rect 19076 15748 19132 15750
rect 19156 15748 19212 15750
rect 19236 15748 19292 15750
rect 18916 14714 18972 14716
rect 18996 14714 19052 14716
rect 19076 14714 19132 14716
rect 19156 14714 19212 14716
rect 19236 14714 19292 14716
rect 18916 14662 18918 14714
rect 18918 14662 18970 14714
rect 18970 14662 18972 14714
rect 18996 14662 19034 14714
rect 19034 14662 19046 14714
rect 19046 14662 19052 14714
rect 19076 14662 19098 14714
rect 19098 14662 19110 14714
rect 19110 14662 19132 14714
rect 19156 14662 19162 14714
rect 19162 14662 19174 14714
rect 19174 14662 19212 14714
rect 19236 14662 19238 14714
rect 19238 14662 19290 14714
rect 19290 14662 19292 14714
rect 18916 14660 18972 14662
rect 18996 14660 19052 14662
rect 19076 14660 19132 14662
rect 19156 14660 19212 14662
rect 19236 14660 19292 14662
rect 19656 16346 19712 16348
rect 19736 16346 19792 16348
rect 19816 16346 19872 16348
rect 19896 16346 19952 16348
rect 19976 16346 20032 16348
rect 19656 16294 19658 16346
rect 19658 16294 19710 16346
rect 19710 16294 19712 16346
rect 19736 16294 19774 16346
rect 19774 16294 19786 16346
rect 19786 16294 19792 16346
rect 19816 16294 19838 16346
rect 19838 16294 19850 16346
rect 19850 16294 19872 16346
rect 19896 16294 19902 16346
rect 19902 16294 19914 16346
rect 19914 16294 19952 16346
rect 19976 16294 19978 16346
rect 19978 16294 20030 16346
rect 20030 16294 20032 16346
rect 19656 16292 19712 16294
rect 19736 16292 19792 16294
rect 19816 16292 19872 16294
rect 19896 16292 19952 16294
rect 19976 16292 20032 16294
rect 19656 15258 19712 15260
rect 19736 15258 19792 15260
rect 19816 15258 19872 15260
rect 19896 15258 19952 15260
rect 19976 15258 20032 15260
rect 19656 15206 19658 15258
rect 19658 15206 19710 15258
rect 19710 15206 19712 15258
rect 19736 15206 19774 15258
rect 19774 15206 19786 15258
rect 19786 15206 19792 15258
rect 19816 15206 19838 15258
rect 19838 15206 19850 15258
rect 19850 15206 19872 15258
rect 19896 15206 19902 15258
rect 19902 15206 19914 15258
rect 19914 15206 19952 15258
rect 19976 15206 19978 15258
rect 19978 15206 20030 15258
rect 20030 15206 20032 15258
rect 19656 15204 19712 15206
rect 19736 15204 19792 15206
rect 19816 15204 19872 15206
rect 19896 15204 19952 15206
rect 19976 15204 20032 15206
rect 18694 14356 18696 14376
rect 18696 14356 18748 14376
rect 18748 14356 18750 14376
rect 18694 14320 18750 14356
rect 18418 13368 18474 13424
rect 19656 14170 19712 14172
rect 19736 14170 19792 14172
rect 19816 14170 19872 14172
rect 19896 14170 19952 14172
rect 19976 14170 20032 14172
rect 19656 14118 19658 14170
rect 19658 14118 19710 14170
rect 19710 14118 19712 14170
rect 19736 14118 19774 14170
rect 19774 14118 19786 14170
rect 19786 14118 19792 14170
rect 19816 14118 19838 14170
rect 19838 14118 19850 14170
rect 19850 14118 19872 14170
rect 19896 14118 19902 14170
rect 19902 14118 19914 14170
rect 19914 14118 19952 14170
rect 19976 14118 19978 14170
rect 19978 14118 20030 14170
rect 20030 14118 20032 14170
rect 19656 14116 19712 14118
rect 19736 14116 19792 14118
rect 19816 14116 19872 14118
rect 19896 14116 19952 14118
rect 19976 14116 20032 14118
rect 18916 13626 18972 13628
rect 18996 13626 19052 13628
rect 19076 13626 19132 13628
rect 19156 13626 19212 13628
rect 19236 13626 19292 13628
rect 18916 13574 18918 13626
rect 18918 13574 18970 13626
rect 18970 13574 18972 13626
rect 18996 13574 19034 13626
rect 19034 13574 19046 13626
rect 19046 13574 19052 13626
rect 19076 13574 19098 13626
rect 19098 13574 19110 13626
rect 19110 13574 19132 13626
rect 19156 13574 19162 13626
rect 19162 13574 19174 13626
rect 19174 13574 19212 13626
rect 19236 13574 19238 13626
rect 19238 13574 19290 13626
rect 19290 13574 19292 13626
rect 18916 13572 18972 13574
rect 18996 13572 19052 13574
rect 19076 13572 19132 13574
rect 19156 13572 19212 13574
rect 19236 13572 19292 13574
rect 18916 12538 18972 12540
rect 18996 12538 19052 12540
rect 19076 12538 19132 12540
rect 19156 12538 19212 12540
rect 19236 12538 19292 12540
rect 18916 12486 18918 12538
rect 18918 12486 18970 12538
rect 18970 12486 18972 12538
rect 18996 12486 19034 12538
rect 19034 12486 19046 12538
rect 19046 12486 19052 12538
rect 19076 12486 19098 12538
rect 19098 12486 19110 12538
rect 19110 12486 19132 12538
rect 19156 12486 19162 12538
rect 19162 12486 19174 12538
rect 19174 12486 19212 12538
rect 19236 12486 19238 12538
rect 19238 12486 19290 12538
rect 19290 12486 19292 12538
rect 18916 12484 18972 12486
rect 18996 12484 19052 12486
rect 19076 12484 19132 12486
rect 19156 12484 19212 12486
rect 19236 12484 19292 12486
rect 19656 13082 19712 13084
rect 19736 13082 19792 13084
rect 19816 13082 19872 13084
rect 19896 13082 19952 13084
rect 19976 13082 20032 13084
rect 19656 13030 19658 13082
rect 19658 13030 19710 13082
rect 19710 13030 19712 13082
rect 19736 13030 19774 13082
rect 19774 13030 19786 13082
rect 19786 13030 19792 13082
rect 19816 13030 19838 13082
rect 19838 13030 19850 13082
rect 19850 13030 19872 13082
rect 19896 13030 19902 13082
rect 19902 13030 19914 13082
rect 19914 13030 19952 13082
rect 19976 13030 19978 13082
rect 19978 13030 20030 13082
rect 20030 13030 20032 13082
rect 19656 13028 19712 13030
rect 19736 13028 19792 13030
rect 19816 13028 19872 13030
rect 19896 13028 19952 13030
rect 19976 13028 20032 13030
rect 18916 11450 18972 11452
rect 18996 11450 19052 11452
rect 19076 11450 19132 11452
rect 19156 11450 19212 11452
rect 19236 11450 19292 11452
rect 18916 11398 18918 11450
rect 18918 11398 18970 11450
rect 18970 11398 18972 11450
rect 18996 11398 19034 11450
rect 19034 11398 19046 11450
rect 19046 11398 19052 11450
rect 19076 11398 19098 11450
rect 19098 11398 19110 11450
rect 19110 11398 19132 11450
rect 19156 11398 19162 11450
rect 19162 11398 19174 11450
rect 19174 11398 19212 11450
rect 19236 11398 19238 11450
rect 19238 11398 19290 11450
rect 19290 11398 19292 11450
rect 18916 11396 18972 11398
rect 18996 11396 19052 11398
rect 19076 11396 19132 11398
rect 19156 11396 19212 11398
rect 19236 11396 19292 11398
rect 18602 10240 18658 10296
rect 18916 10362 18972 10364
rect 18996 10362 19052 10364
rect 19076 10362 19132 10364
rect 19156 10362 19212 10364
rect 19236 10362 19292 10364
rect 18916 10310 18918 10362
rect 18918 10310 18970 10362
rect 18970 10310 18972 10362
rect 18996 10310 19034 10362
rect 19034 10310 19046 10362
rect 19046 10310 19052 10362
rect 19076 10310 19098 10362
rect 19098 10310 19110 10362
rect 19110 10310 19132 10362
rect 19156 10310 19162 10362
rect 19162 10310 19174 10362
rect 19174 10310 19212 10362
rect 19236 10310 19238 10362
rect 19238 10310 19290 10362
rect 19290 10310 19292 10362
rect 18916 10308 18972 10310
rect 18996 10308 19052 10310
rect 19076 10308 19132 10310
rect 19156 10308 19212 10310
rect 19236 10308 19292 10310
rect 19656 11994 19712 11996
rect 19736 11994 19792 11996
rect 19816 11994 19872 11996
rect 19896 11994 19952 11996
rect 19976 11994 20032 11996
rect 19656 11942 19658 11994
rect 19658 11942 19710 11994
rect 19710 11942 19712 11994
rect 19736 11942 19774 11994
rect 19774 11942 19786 11994
rect 19786 11942 19792 11994
rect 19816 11942 19838 11994
rect 19838 11942 19850 11994
rect 19850 11942 19872 11994
rect 19896 11942 19902 11994
rect 19902 11942 19914 11994
rect 19914 11942 19952 11994
rect 19976 11942 19978 11994
rect 19978 11942 20030 11994
rect 20030 11942 20032 11994
rect 19656 11940 19712 11942
rect 19736 11940 19792 11942
rect 19816 11940 19872 11942
rect 19896 11940 19952 11942
rect 19976 11940 20032 11942
rect 19656 10906 19712 10908
rect 19736 10906 19792 10908
rect 19816 10906 19872 10908
rect 19896 10906 19952 10908
rect 19976 10906 20032 10908
rect 19656 10854 19658 10906
rect 19658 10854 19710 10906
rect 19710 10854 19712 10906
rect 19736 10854 19774 10906
rect 19774 10854 19786 10906
rect 19786 10854 19792 10906
rect 19816 10854 19838 10906
rect 19838 10854 19850 10906
rect 19850 10854 19872 10906
rect 19896 10854 19902 10906
rect 19902 10854 19914 10906
rect 19914 10854 19952 10906
rect 19976 10854 19978 10906
rect 19978 10854 20030 10906
rect 20030 10854 20032 10906
rect 19656 10852 19712 10854
rect 19736 10852 19792 10854
rect 19816 10852 19872 10854
rect 19896 10852 19952 10854
rect 19976 10852 20032 10854
rect 20718 22072 20774 22128
rect 22916 27770 22972 27772
rect 22996 27770 23052 27772
rect 23076 27770 23132 27772
rect 23156 27770 23212 27772
rect 23236 27770 23292 27772
rect 22916 27718 22918 27770
rect 22918 27718 22970 27770
rect 22970 27718 22972 27770
rect 22996 27718 23034 27770
rect 23034 27718 23046 27770
rect 23046 27718 23052 27770
rect 23076 27718 23098 27770
rect 23098 27718 23110 27770
rect 23110 27718 23132 27770
rect 23156 27718 23162 27770
rect 23162 27718 23174 27770
rect 23174 27718 23212 27770
rect 23236 27718 23238 27770
rect 23238 27718 23290 27770
rect 23290 27718 23292 27770
rect 22916 27716 22972 27718
rect 22996 27716 23052 27718
rect 23076 27716 23132 27718
rect 23156 27716 23212 27718
rect 23236 27716 23292 27718
rect 23656 27226 23712 27228
rect 23736 27226 23792 27228
rect 23816 27226 23872 27228
rect 23896 27226 23952 27228
rect 23976 27226 24032 27228
rect 23656 27174 23658 27226
rect 23658 27174 23710 27226
rect 23710 27174 23712 27226
rect 23736 27174 23774 27226
rect 23774 27174 23786 27226
rect 23786 27174 23792 27226
rect 23816 27174 23838 27226
rect 23838 27174 23850 27226
rect 23850 27174 23872 27226
rect 23896 27174 23902 27226
rect 23902 27174 23914 27226
rect 23914 27174 23952 27226
rect 23976 27174 23978 27226
rect 23978 27174 24030 27226
rect 24030 27174 24032 27226
rect 23656 27172 23712 27174
rect 23736 27172 23792 27174
rect 23816 27172 23872 27174
rect 23896 27172 23952 27174
rect 23976 27172 24032 27174
rect 22916 26682 22972 26684
rect 22996 26682 23052 26684
rect 23076 26682 23132 26684
rect 23156 26682 23212 26684
rect 23236 26682 23292 26684
rect 22916 26630 22918 26682
rect 22918 26630 22970 26682
rect 22970 26630 22972 26682
rect 22996 26630 23034 26682
rect 23034 26630 23046 26682
rect 23046 26630 23052 26682
rect 23076 26630 23098 26682
rect 23098 26630 23110 26682
rect 23110 26630 23132 26682
rect 23156 26630 23162 26682
rect 23162 26630 23174 26682
rect 23174 26630 23212 26682
rect 23236 26630 23238 26682
rect 23238 26630 23290 26682
rect 23290 26630 23292 26682
rect 22916 26628 22972 26630
rect 22996 26628 23052 26630
rect 23076 26628 23132 26630
rect 23156 26628 23212 26630
rect 23236 26628 23292 26630
rect 23656 26138 23712 26140
rect 23736 26138 23792 26140
rect 23816 26138 23872 26140
rect 23896 26138 23952 26140
rect 23976 26138 24032 26140
rect 23656 26086 23658 26138
rect 23658 26086 23710 26138
rect 23710 26086 23712 26138
rect 23736 26086 23774 26138
rect 23774 26086 23786 26138
rect 23786 26086 23792 26138
rect 23816 26086 23838 26138
rect 23838 26086 23850 26138
rect 23850 26086 23872 26138
rect 23896 26086 23902 26138
rect 23902 26086 23914 26138
rect 23914 26086 23952 26138
rect 23976 26086 23978 26138
rect 23978 26086 24030 26138
rect 24030 26086 24032 26138
rect 23656 26084 23712 26086
rect 23736 26084 23792 26086
rect 23816 26084 23872 26086
rect 23896 26084 23952 26086
rect 23976 26084 24032 26086
rect 22916 25594 22972 25596
rect 22996 25594 23052 25596
rect 23076 25594 23132 25596
rect 23156 25594 23212 25596
rect 23236 25594 23292 25596
rect 22916 25542 22918 25594
rect 22918 25542 22970 25594
rect 22970 25542 22972 25594
rect 22996 25542 23034 25594
rect 23034 25542 23046 25594
rect 23046 25542 23052 25594
rect 23076 25542 23098 25594
rect 23098 25542 23110 25594
rect 23110 25542 23132 25594
rect 23156 25542 23162 25594
rect 23162 25542 23174 25594
rect 23174 25542 23212 25594
rect 23236 25542 23238 25594
rect 23238 25542 23290 25594
rect 23290 25542 23292 25594
rect 22916 25540 22972 25542
rect 22996 25540 23052 25542
rect 23076 25540 23132 25542
rect 23156 25540 23212 25542
rect 23236 25540 23292 25542
rect 22916 24506 22972 24508
rect 22996 24506 23052 24508
rect 23076 24506 23132 24508
rect 23156 24506 23212 24508
rect 23236 24506 23292 24508
rect 22916 24454 22918 24506
rect 22918 24454 22970 24506
rect 22970 24454 22972 24506
rect 22996 24454 23034 24506
rect 23034 24454 23046 24506
rect 23046 24454 23052 24506
rect 23076 24454 23098 24506
rect 23098 24454 23110 24506
rect 23110 24454 23132 24506
rect 23156 24454 23162 24506
rect 23162 24454 23174 24506
rect 23174 24454 23212 24506
rect 23236 24454 23238 24506
rect 23238 24454 23290 24506
rect 23290 24454 23292 24506
rect 22916 24452 22972 24454
rect 22996 24452 23052 24454
rect 23076 24452 23132 24454
rect 23156 24452 23212 24454
rect 23236 24452 23292 24454
rect 22916 23418 22972 23420
rect 22996 23418 23052 23420
rect 23076 23418 23132 23420
rect 23156 23418 23212 23420
rect 23236 23418 23292 23420
rect 22916 23366 22918 23418
rect 22918 23366 22970 23418
rect 22970 23366 22972 23418
rect 22996 23366 23034 23418
rect 23034 23366 23046 23418
rect 23046 23366 23052 23418
rect 23076 23366 23098 23418
rect 23098 23366 23110 23418
rect 23110 23366 23132 23418
rect 23156 23366 23162 23418
rect 23162 23366 23174 23418
rect 23174 23366 23212 23418
rect 23236 23366 23238 23418
rect 23238 23366 23290 23418
rect 23290 23366 23292 23418
rect 22916 23364 22972 23366
rect 22996 23364 23052 23366
rect 23076 23364 23132 23366
rect 23156 23364 23212 23366
rect 23236 23364 23292 23366
rect 23656 25050 23712 25052
rect 23736 25050 23792 25052
rect 23816 25050 23872 25052
rect 23896 25050 23952 25052
rect 23976 25050 24032 25052
rect 23656 24998 23658 25050
rect 23658 24998 23710 25050
rect 23710 24998 23712 25050
rect 23736 24998 23774 25050
rect 23774 24998 23786 25050
rect 23786 24998 23792 25050
rect 23816 24998 23838 25050
rect 23838 24998 23850 25050
rect 23850 24998 23872 25050
rect 23896 24998 23902 25050
rect 23902 24998 23914 25050
rect 23914 24998 23952 25050
rect 23976 24998 23978 25050
rect 23978 24998 24030 25050
rect 24030 24998 24032 25050
rect 23656 24996 23712 24998
rect 23736 24996 23792 24998
rect 23816 24996 23872 24998
rect 23896 24996 23952 24998
rect 23976 24996 24032 24998
rect 24490 24928 24546 24984
rect 23656 23962 23712 23964
rect 23736 23962 23792 23964
rect 23816 23962 23872 23964
rect 23896 23962 23952 23964
rect 23976 23962 24032 23964
rect 23656 23910 23658 23962
rect 23658 23910 23710 23962
rect 23710 23910 23712 23962
rect 23736 23910 23774 23962
rect 23774 23910 23786 23962
rect 23786 23910 23792 23962
rect 23816 23910 23838 23962
rect 23838 23910 23850 23962
rect 23850 23910 23872 23962
rect 23896 23910 23902 23962
rect 23902 23910 23914 23962
rect 23914 23910 23952 23962
rect 23976 23910 23978 23962
rect 23978 23910 24030 23962
rect 24030 23910 24032 23962
rect 23656 23908 23712 23910
rect 23736 23908 23792 23910
rect 23816 23908 23872 23910
rect 23896 23908 23952 23910
rect 23976 23908 24032 23910
rect 23656 22874 23712 22876
rect 23736 22874 23792 22876
rect 23816 22874 23872 22876
rect 23896 22874 23952 22876
rect 23976 22874 24032 22876
rect 23656 22822 23658 22874
rect 23658 22822 23710 22874
rect 23710 22822 23712 22874
rect 23736 22822 23774 22874
rect 23774 22822 23786 22874
rect 23786 22822 23792 22874
rect 23816 22822 23838 22874
rect 23838 22822 23850 22874
rect 23850 22822 23872 22874
rect 23896 22822 23902 22874
rect 23902 22822 23914 22874
rect 23914 22822 23952 22874
rect 23976 22822 23978 22874
rect 23978 22822 24030 22874
rect 24030 22822 24032 22874
rect 23656 22820 23712 22822
rect 23736 22820 23792 22822
rect 23816 22820 23872 22822
rect 23896 22820 23952 22822
rect 23976 22820 24032 22822
rect 22916 22330 22972 22332
rect 22996 22330 23052 22332
rect 23076 22330 23132 22332
rect 23156 22330 23212 22332
rect 23236 22330 23292 22332
rect 22916 22278 22918 22330
rect 22918 22278 22970 22330
rect 22970 22278 22972 22330
rect 22996 22278 23034 22330
rect 23034 22278 23046 22330
rect 23046 22278 23052 22330
rect 23076 22278 23098 22330
rect 23098 22278 23110 22330
rect 23110 22278 23132 22330
rect 23156 22278 23162 22330
rect 23162 22278 23174 22330
rect 23174 22278 23212 22330
rect 23236 22278 23238 22330
rect 23238 22278 23290 22330
rect 23290 22278 23292 22330
rect 22916 22276 22972 22278
rect 22996 22276 23052 22278
rect 23076 22276 23132 22278
rect 23156 22276 23212 22278
rect 23236 22276 23292 22278
rect 22916 21242 22972 21244
rect 22996 21242 23052 21244
rect 23076 21242 23132 21244
rect 23156 21242 23212 21244
rect 23236 21242 23292 21244
rect 22916 21190 22918 21242
rect 22918 21190 22970 21242
rect 22970 21190 22972 21242
rect 22996 21190 23034 21242
rect 23034 21190 23046 21242
rect 23046 21190 23052 21242
rect 23076 21190 23098 21242
rect 23098 21190 23110 21242
rect 23110 21190 23132 21242
rect 23156 21190 23162 21242
rect 23162 21190 23174 21242
rect 23174 21190 23212 21242
rect 23236 21190 23238 21242
rect 23238 21190 23290 21242
rect 23290 21190 23292 21242
rect 22916 21188 22972 21190
rect 22996 21188 23052 21190
rect 23076 21188 23132 21190
rect 23156 21188 23212 21190
rect 23236 21188 23292 21190
rect 23656 21786 23712 21788
rect 23736 21786 23792 21788
rect 23816 21786 23872 21788
rect 23896 21786 23952 21788
rect 23976 21786 24032 21788
rect 23656 21734 23658 21786
rect 23658 21734 23710 21786
rect 23710 21734 23712 21786
rect 23736 21734 23774 21786
rect 23774 21734 23786 21786
rect 23786 21734 23792 21786
rect 23816 21734 23838 21786
rect 23838 21734 23850 21786
rect 23850 21734 23872 21786
rect 23896 21734 23902 21786
rect 23902 21734 23914 21786
rect 23914 21734 23952 21786
rect 23976 21734 23978 21786
rect 23978 21734 24030 21786
rect 24030 21734 24032 21786
rect 23656 21732 23712 21734
rect 23736 21732 23792 21734
rect 23816 21732 23872 21734
rect 23896 21732 23952 21734
rect 23976 21732 24032 21734
rect 22916 20154 22972 20156
rect 22996 20154 23052 20156
rect 23076 20154 23132 20156
rect 23156 20154 23212 20156
rect 23236 20154 23292 20156
rect 22916 20102 22918 20154
rect 22918 20102 22970 20154
rect 22970 20102 22972 20154
rect 22996 20102 23034 20154
rect 23034 20102 23046 20154
rect 23046 20102 23052 20154
rect 23076 20102 23098 20154
rect 23098 20102 23110 20154
rect 23110 20102 23132 20154
rect 23156 20102 23162 20154
rect 23162 20102 23174 20154
rect 23174 20102 23212 20154
rect 23236 20102 23238 20154
rect 23238 20102 23290 20154
rect 23290 20102 23292 20154
rect 22916 20100 22972 20102
rect 22996 20100 23052 20102
rect 23076 20100 23132 20102
rect 23156 20100 23212 20102
rect 23236 20100 23292 20102
rect 23656 20698 23712 20700
rect 23736 20698 23792 20700
rect 23816 20698 23872 20700
rect 23896 20698 23952 20700
rect 23976 20698 24032 20700
rect 23656 20646 23658 20698
rect 23658 20646 23710 20698
rect 23710 20646 23712 20698
rect 23736 20646 23774 20698
rect 23774 20646 23786 20698
rect 23786 20646 23792 20698
rect 23816 20646 23838 20698
rect 23838 20646 23850 20698
rect 23850 20646 23872 20698
rect 23896 20646 23902 20698
rect 23902 20646 23914 20698
rect 23914 20646 23952 20698
rect 23976 20646 23978 20698
rect 23978 20646 24030 20698
rect 24030 20646 24032 20698
rect 23656 20644 23712 20646
rect 23736 20644 23792 20646
rect 23816 20644 23872 20646
rect 23896 20644 23952 20646
rect 23976 20644 24032 20646
rect 19656 9818 19712 9820
rect 19736 9818 19792 9820
rect 19816 9818 19872 9820
rect 19896 9818 19952 9820
rect 19976 9818 20032 9820
rect 19656 9766 19658 9818
rect 19658 9766 19710 9818
rect 19710 9766 19712 9818
rect 19736 9766 19774 9818
rect 19774 9766 19786 9818
rect 19786 9766 19792 9818
rect 19816 9766 19838 9818
rect 19838 9766 19850 9818
rect 19850 9766 19872 9818
rect 19896 9766 19902 9818
rect 19902 9766 19914 9818
rect 19914 9766 19952 9818
rect 19976 9766 19978 9818
rect 19978 9766 20030 9818
rect 20030 9766 20032 9818
rect 19656 9764 19712 9766
rect 19736 9764 19792 9766
rect 19816 9764 19872 9766
rect 19896 9764 19952 9766
rect 19976 9764 20032 9766
rect 10916 2746 10972 2748
rect 10996 2746 11052 2748
rect 11076 2746 11132 2748
rect 11156 2746 11212 2748
rect 11236 2746 11292 2748
rect 10916 2694 10918 2746
rect 10918 2694 10970 2746
rect 10970 2694 10972 2746
rect 10996 2694 11034 2746
rect 11034 2694 11046 2746
rect 11046 2694 11052 2746
rect 11076 2694 11098 2746
rect 11098 2694 11110 2746
rect 11110 2694 11132 2746
rect 11156 2694 11162 2746
rect 11162 2694 11174 2746
rect 11174 2694 11212 2746
rect 11236 2694 11238 2746
rect 11238 2694 11290 2746
rect 11290 2694 11292 2746
rect 10916 2692 10972 2694
rect 10996 2692 11052 2694
rect 11076 2692 11132 2694
rect 11156 2692 11212 2694
rect 11236 2692 11292 2694
rect 14916 2746 14972 2748
rect 14996 2746 15052 2748
rect 15076 2746 15132 2748
rect 15156 2746 15212 2748
rect 15236 2746 15292 2748
rect 14916 2694 14918 2746
rect 14918 2694 14970 2746
rect 14970 2694 14972 2746
rect 14996 2694 15034 2746
rect 15034 2694 15046 2746
rect 15046 2694 15052 2746
rect 15076 2694 15098 2746
rect 15098 2694 15110 2746
rect 15110 2694 15132 2746
rect 15156 2694 15162 2746
rect 15162 2694 15174 2746
rect 15174 2694 15212 2746
rect 15236 2694 15238 2746
rect 15238 2694 15290 2746
rect 15290 2694 15292 2746
rect 14916 2692 14972 2694
rect 14996 2692 15052 2694
rect 15076 2692 15132 2694
rect 15156 2692 15212 2694
rect 15236 2692 15292 2694
rect 18916 9274 18972 9276
rect 18996 9274 19052 9276
rect 19076 9274 19132 9276
rect 19156 9274 19212 9276
rect 19236 9274 19292 9276
rect 18916 9222 18918 9274
rect 18918 9222 18970 9274
rect 18970 9222 18972 9274
rect 18996 9222 19034 9274
rect 19034 9222 19046 9274
rect 19046 9222 19052 9274
rect 19076 9222 19098 9274
rect 19098 9222 19110 9274
rect 19110 9222 19132 9274
rect 19156 9222 19162 9274
rect 19162 9222 19174 9274
rect 19174 9222 19212 9274
rect 19236 9222 19238 9274
rect 19238 9222 19290 9274
rect 19290 9222 19292 9274
rect 18916 9220 18972 9222
rect 18996 9220 19052 9222
rect 19076 9220 19132 9222
rect 19156 9220 19212 9222
rect 19236 9220 19292 9222
rect 18916 8186 18972 8188
rect 18996 8186 19052 8188
rect 19076 8186 19132 8188
rect 19156 8186 19212 8188
rect 19236 8186 19292 8188
rect 18916 8134 18918 8186
rect 18918 8134 18970 8186
rect 18970 8134 18972 8186
rect 18996 8134 19034 8186
rect 19034 8134 19046 8186
rect 19046 8134 19052 8186
rect 19076 8134 19098 8186
rect 19098 8134 19110 8186
rect 19110 8134 19132 8186
rect 19156 8134 19162 8186
rect 19162 8134 19174 8186
rect 19174 8134 19212 8186
rect 19236 8134 19238 8186
rect 19238 8134 19290 8186
rect 19290 8134 19292 8186
rect 18916 8132 18972 8134
rect 18996 8132 19052 8134
rect 19076 8132 19132 8134
rect 19156 8132 19212 8134
rect 19236 8132 19292 8134
rect 18916 7098 18972 7100
rect 18996 7098 19052 7100
rect 19076 7098 19132 7100
rect 19156 7098 19212 7100
rect 19236 7098 19292 7100
rect 18916 7046 18918 7098
rect 18918 7046 18970 7098
rect 18970 7046 18972 7098
rect 18996 7046 19034 7098
rect 19034 7046 19046 7098
rect 19046 7046 19052 7098
rect 19076 7046 19098 7098
rect 19098 7046 19110 7098
rect 19110 7046 19132 7098
rect 19156 7046 19162 7098
rect 19162 7046 19174 7098
rect 19174 7046 19212 7098
rect 19236 7046 19238 7098
rect 19238 7046 19290 7098
rect 19290 7046 19292 7098
rect 18916 7044 18972 7046
rect 18996 7044 19052 7046
rect 19076 7044 19132 7046
rect 19156 7044 19212 7046
rect 19236 7044 19292 7046
rect 19656 8730 19712 8732
rect 19736 8730 19792 8732
rect 19816 8730 19872 8732
rect 19896 8730 19952 8732
rect 19976 8730 20032 8732
rect 19656 8678 19658 8730
rect 19658 8678 19710 8730
rect 19710 8678 19712 8730
rect 19736 8678 19774 8730
rect 19774 8678 19786 8730
rect 19786 8678 19792 8730
rect 19816 8678 19838 8730
rect 19838 8678 19850 8730
rect 19850 8678 19872 8730
rect 19896 8678 19902 8730
rect 19902 8678 19914 8730
rect 19914 8678 19952 8730
rect 19976 8678 19978 8730
rect 19978 8678 20030 8730
rect 20030 8678 20032 8730
rect 19656 8676 19712 8678
rect 19736 8676 19792 8678
rect 19816 8676 19872 8678
rect 19896 8676 19952 8678
rect 19976 8676 20032 8678
rect 19706 7964 19708 7984
rect 19708 7964 19760 7984
rect 19760 7964 19762 7984
rect 19706 7928 19762 7964
rect 19656 7642 19712 7644
rect 19736 7642 19792 7644
rect 19816 7642 19872 7644
rect 19896 7642 19952 7644
rect 19976 7642 20032 7644
rect 19656 7590 19658 7642
rect 19658 7590 19710 7642
rect 19710 7590 19712 7642
rect 19736 7590 19774 7642
rect 19774 7590 19786 7642
rect 19786 7590 19792 7642
rect 19816 7590 19838 7642
rect 19838 7590 19850 7642
rect 19850 7590 19872 7642
rect 19896 7590 19902 7642
rect 19902 7590 19914 7642
rect 19914 7590 19952 7642
rect 19976 7590 19978 7642
rect 19978 7590 20030 7642
rect 20030 7590 20032 7642
rect 19656 7588 19712 7590
rect 19736 7588 19792 7590
rect 19816 7588 19872 7590
rect 19896 7588 19952 7590
rect 19976 7588 20032 7590
rect 18916 6010 18972 6012
rect 18996 6010 19052 6012
rect 19076 6010 19132 6012
rect 19156 6010 19212 6012
rect 19236 6010 19292 6012
rect 18916 5958 18918 6010
rect 18918 5958 18970 6010
rect 18970 5958 18972 6010
rect 18996 5958 19034 6010
rect 19034 5958 19046 6010
rect 19046 5958 19052 6010
rect 19076 5958 19098 6010
rect 19098 5958 19110 6010
rect 19110 5958 19132 6010
rect 19156 5958 19162 6010
rect 19162 5958 19174 6010
rect 19174 5958 19212 6010
rect 19236 5958 19238 6010
rect 19238 5958 19290 6010
rect 19290 5958 19292 6010
rect 18916 5956 18972 5958
rect 18996 5956 19052 5958
rect 19076 5956 19132 5958
rect 19156 5956 19212 5958
rect 19236 5956 19292 5958
rect 19656 6554 19712 6556
rect 19736 6554 19792 6556
rect 19816 6554 19872 6556
rect 19896 6554 19952 6556
rect 19976 6554 20032 6556
rect 19656 6502 19658 6554
rect 19658 6502 19710 6554
rect 19710 6502 19712 6554
rect 19736 6502 19774 6554
rect 19774 6502 19786 6554
rect 19786 6502 19792 6554
rect 19816 6502 19838 6554
rect 19838 6502 19850 6554
rect 19850 6502 19872 6554
rect 19896 6502 19902 6554
rect 19902 6502 19914 6554
rect 19914 6502 19952 6554
rect 19976 6502 19978 6554
rect 19978 6502 20030 6554
rect 20030 6502 20032 6554
rect 19656 6500 19712 6502
rect 19736 6500 19792 6502
rect 19816 6500 19872 6502
rect 19896 6500 19952 6502
rect 19976 6500 20032 6502
rect 18916 4922 18972 4924
rect 18996 4922 19052 4924
rect 19076 4922 19132 4924
rect 19156 4922 19212 4924
rect 19236 4922 19292 4924
rect 18916 4870 18918 4922
rect 18918 4870 18970 4922
rect 18970 4870 18972 4922
rect 18996 4870 19034 4922
rect 19034 4870 19046 4922
rect 19046 4870 19052 4922
rect 19076 4870 19098 4922
rect 19098 4870 19110 4922
rect 19110 4870 19132 4922
rect 19156 4870 19162 4922
rect 19162 4870 19174 4922
rect 19174 4870 19212 4922
rect 19236 4870 19238 4922
rect 19238 4870 19290 4922
rect 19290 4870 19292 4922
rect 18916 4868 18972 4870
rect 18996 4868 19052 4870
rect 19076 4868 19132 4870
rect 19156 4868 19212 4870
rect 19236 4868 19292 4870
rect 18916 3834 18972 3836
rect 18996 3834 19052 3836
rect 19076 3834 19132 3836
rect 19156 3834 19212 3836
rect 19236 3834 19292 3836
rect 18916 3782 18918 3834
rect 18918 3782 18970 3834
rect 18970 3782 18972 3834
rect 18996 3782 19034 3834
rect 19034 3782 19046 3834
rect 19046 3782 19052 3834
rect 19076 3782 19098 3834
rect 19098 3782 19110 3834
rect 19110 3782 19132 3834
rect 19156 3782 19162 3834
rect 19162 3782 19174 3834
rect 19174 3782 19212 3834
rect 19236 3782 19238 3834
rect 19238 3782 19290 3834
rect 19290 3782 19292 3834
rect 18916 3780 18972 3782
rect 18996 3780 19052 3782
rect 19076 3780 19132 3782
rect 19156 3780 19212 3782
rect 19236 3780 19292 3782
rect 18916 2746 18972 2748
rect 18996 2746 19052 2748
rect 19076 2746 19132 2748
rect 19156 2746 19212 2748
rect 19236 2746 19292 2748
rect 18916 2694 18918 2746
rect 18918 2694 18970 2746
rect 18970 2694 18972 2746
rect 18996 2694 19034 2746
rect 19034 2694 19046 2746
rect 19046 2694 19052 2746
rect 19076 2694 19098 2746
rect 19098 2694 19110 2746
rect 19110 2694 19132 2746
rect 19156 2694 19162 2746
rect 19162 2694 19174 2746
rect 19174 2694 19212 2746
rect 19236 2694 19238 2746
rect 19238 2694 19290 2746
rect 19290 2694 19292 2746
rect 18916 2692 18972 2694
rect 18996 2692 19052 2694
rect 19076 2692 19132 2694
rect 19156 2692 19212 2694
rect 19236 2692 19292 2694
rect 3656 2202 3712 2204
rect 3736 2202 3792 2204
rect 3816 2202 3872 2204
rect 3896 2202 3952 2204
rect 3976 2202 4032 2204
rect 3656 2150 3658 2202
rect 3658 2150 3710 2202
rect 3710 2150 3712 2202
rect 3736 2150 3774 2202
rect 3774 2150 3786 2202
rect 3786 2150 3792 2202
rect 3816 2150 3838 2202
rect 3838 2150 3850 2202
rect 3850 2150 3872 2202
rect 3896 2150 3902 2202
rect 3902 2150 3914 2202
rect 3914 2150 3952 2202
rect 3976 2150 3978 2202
rect 3978 2150 4030 2202
rect 4030 2150 4032 2202
rect 3656 2148 3712 2150
rect 3736 2148 3792 2150
rect 3816 2148 3872 2150
rect 3896 2148 3952 2150
rect 3976 2148 4032 2150
rect 7656 2202 7712 2204
rect 7736 2202 7792 2204
rect 7816 2202 7872 2204
rect 7896 2202 7952 2204
rect 7976 2202 8032 2204
rect 7656 2150 7658 2202
rect 7658 2150 7710 2202
rect 7710 2150 7712 2202
rect 7736 2150 7774 2202
rect 7774 2150 7786 2202
rect 7786 2150 7792 2202
rect 7816 2150 7838 2202
rect 7838 2150 7850 2202
rect 7850 2150 7872 2202
rect 7896 2150 7902 2202
rect 7902 2150 7914 2202
rect 7914 2150 7952 2202
rect 7976 2150 7978 2202
rect 7978 2150 8030 2202
rect 8030 2150 8032 2202
rect 7656 2148 7712 2150
rect 7736 2148 7792 2150
rect 7816 2148 7872 2150
rect 7896 2148 7952 2150
rect 7976 2148 8032 2150
rect 11656 2202 11712 2204
rect 11736 2202 11792 2204
rect 11816 2202 11872 2204
rect 11896 2202 11952 2204
rect 11976 2202 12032 2204
rect 11656 2150 11658 2202
rect 11658 2150 11710 2202
rect 11710 2150 11712 2202
rect 11736 2150 11774 2202
rect 11774 2150 11786 2202
rect 11786 2150 11792 2202
rect 11816 2150 11838 2202
rect 11838 2150 11850 2202
rect 11850 2150 11872 2202
rect 11896 2150 11902 2202
rect 11902 2150 11914 2202
rect 11914 2150 11952 2202
rect 11976 2150 11978 2202
rect 11978 2150 12030 2202
rect 12030 2150 12032 2202
rect 11656 2148 11712 2150
rect 11736 2148 11792 2150
rect 11816 2148 11872 2150
rect 11896 2148 11952 2150
rect 11976 2148 12032 2150
rect 15656 2202 15712 2204
rect 15736 2202 15792 2204
rect 15816 2202 15872 2204
rect 15896 2202 15952 2204
rect 15976 2202 16032 2204
rect 15656 2150 15658 2202
rect 15658 2150 15710 2202
rect 15710 2150 15712 2202
rect 15736 2150 15774 2202
rect 15774 2150 15786 2202
rect 15786 2150 15792 2202
rect 15816 2150 15838 2202
rect 15838 2150 15850 2202
rect 15850 2150 15872 2202
rect 15896 2150 15902 2202
rect 15902 2150 15914 2202
rect 15914 2150 15952 2202
rect 15976 2150 15978 2202
rect 15978 2150 16030 2202
rect 16030 2150 16032 2202
rect 15656 2148 15712 2150
rect 15736 2148 15792 2150
rect 15816 2148 15872 2150
rect 15896 2148 15952 2150
rect 15976 2148 16032 2150
rect 21822 16124 21824 16144
rect 21824 16124 21876 16144
rect 21876 16124 21878 16144
rect 21822 16088 21878 16124
rect 22916 19066 22972 19068
rect 22996 19066 23052 19068
rect 23076 19066 23132 19068
rect 23156 19066 23212 19068
rect 23236 19066 23292 19068
rect 22916 19014 22918 19066
rect 22918 19014 22970 19066
rect 22970 19014 22972 19066
rect 22996 19014 23034 19066
rect 23034 19014 23046 19066
rect 23046 19014 23052 19066
rect 23076 19014 23098 19066
rect 23098 19014 23110 19066
rect 23110 19014 23132 19066
rect 23156 19014 23162 19066
rect 23162 19014 23174 19066
rect 23174 19014 23212 19066
rect 23236 19014 23238 19066
rect 23238 19014 23290 19066
rect 23290 19014 23292 19066
rect 22916 19012 22972 19014
rect 22996 19012 23052 19014
rect 23076 19012 23132 19014
rect 23156 19012 23212 19014
rect 23236 19012 23292 19014
rect 22916 17978 22972 17980
rect 22996 17978 23052 17980
rect 23076 17978 23132 17980
rect 23156 17978 23212 17980
rect 23236 17978 23292 17980
rect 22916 17926 22918 17978
rect 22918 17926 22970 17978
rect 22970 17926 22972 17978
rect 22996 17926 23034 17978
rect 23034 17926 23046 17978
rect 23046 17926 23052 17978
rect 23076 17926 23098 17978
rect 23098 17926 23110 17978
rect 23110 17926 23132 17978
rect 23156 17926 23162 17978
rect 23162 17926 23174 17978
rect 23174 17926 23212 17978
rect 23236 17926 23238 17978
rect 23238 17926 23290 17978
rect 23290 17926 23292 17978
rect 22916 17924 22972 17926
rect 22996 17924 23052 17926
rect 23076 17924 23132 17926
rect 23156 17924 23212 17926
rect 23236 17924 23292 17926
rect 22916 16890 22972 16892
rect 22996 16890 23052 16892
rect 23076 16890 23132 16892
rect 23156 16890 23212 16892
rect 23236 16890 23292 16892
rect 22916 16838 22918 16890
rect 22918 16838 22970 16890
rect 22970 16838 22972 16890
rect 22996 16838 23034 16890
rect 23034 16838 23046 16890
rect 23046 16838 23052 16890
rect 23076 16838 23098 16890
rect 23098 16838 23110 16890
rect 23110 16838 23132 16890
rect 23156 16838 23162 16890
rect 23162 16838 23174 16890
rect 23174 16838 23212 16890
rect 23236 16838 23238 16890
rect 23238 16838 23290 16890
rect 23290 16838 23292 16890
rect 22916 16836 22972 16838
rect 22996 16836 23052 16838
rect 23076 16836 23132 16838
rect 23156 16836 23212 16838
rect 23236 16836 23292 16838
rect 22916 15802 22972 15804
rect 22996 15802 23052 15804
rect 23076 15802 23132 15804
rect 23156 15802 23212 15804
rect 23236 15802 23292 15804
rect 22916 15750 22918 15802
rect 22918 15750 22970 15802
rect 22970 15750 22972 15802
rect 22996 15750 23034 15802
rect 23034 15750 23046 15802
rect 23046 15750 23052 15802
rect 23076 15750 23098 15802
rect 23098 15750 23110 15802
rect 23110 15750 23132 15802
rect 23156 15750 23162 15802
rect 23162 15750 23174 15802
rect 23174 15750 23212 15802
rect 23236 15750 23238 15802
rect 23238 15750 23290 15802
rect 23290 15750 23292 15802
rect 22916 15748 22972 15750
rect 22996 15748 23052 15750
rect 23076 15748 23132 15750
rect 23156 15748 23212 15750
rect 23236 15748 23292 15750
rect 22916 14714 22972 14716
rect 22996 14714 23052 14716
rect 23076 14714 23132 14716
rect 23156 14714 23212 14716
rect 23236 14714 23292 14716
rect 22916 14662 22918 14714
rect 22918 14662 22970 14714
rect 22970 14662 22972 14714
rect 22996 14662 23034 14714
rect 23034 14662 23046 14714
rect 23046 14662 23052 14714
rect 23076 14662 23098 14714
rect 23098 14662 23110 14714
rect 23110 14662 23132 14714
rect 23156 14662 23162 14714
rect 23162 14662 23174 14714
rect 23174 14662 23212 14714
rect 23236 14662 23238 14714
rect 23238 14662 23290 14714
rect 23290 14662 23292 14714
rect 22916 14660 22972 14662
rect 22996 14660 23052 14662
rect 23076 14660 23132 14662
rect 23156 14660 23212 14662
rect 23236 14660 23292 14662
rect 22916 13626 22972 13628
rect 22996 13626 23052 13628
rect 23076 13626 23132 13628
rect 23156 13626 23212 13628
rect 23236 13626 23292 13628
rect 22916 13574 22918 13626
rect 22918 13574 22970 13626
rect 22970 13574 22972 13626
rect 22996 13574 23034 13626
rect 23034 13574 23046 13626
rect 23046 13574 23052 13626
rect 23076 13574 23098 13626
rect 23098 13574 23110 13626
rect 23110 13574 23132 13626
rect 23156 13574 23162 13626
rect 23162 13574 23174 13626
rect 23174 13574 23212 13626
rect 23236 13574 23238 13626
rect 23238 13574 23290 13626
rect 23290 13574 23292 13626
rect 22916 13572 22972 13574
rect 22996 13572 23052 13574
rect 23076 13572 23132 13574
rect 23156 13572 23212 13574
rect 23236 13572 23292 13574
rect 22916 12538 22972 12540
rect 22996 12538 23052 12540
rect 23076 12538 23132 12540
rect 23156 12538 23212 12540
rect 23236 12538 23292 12540
rect 22916 12486 22918 12538
rect 22918 12486 22970 12538
rect 22970 12486 22972 12538
rect 22996 12486 23034 12538
rect 23034 12486 23046 12538
rect 23046 12486 23052 12538
rect 23076 12486 23098 12538
rect 23098 12486 23110 12538
rect 23110 12486 23132 12538
rect 23156 12486 23162 12538
rect 23162 12486 23174 12538
rect 23174 12486 23212 12538
rect 23236 12486 23238 12538
rect 23238 12486 23290 12538
rect 23290 12486 23292 12538
rect 22916 12484 22972 12486
rect 22996 12484 23052 12486
rect 23076 12484 23132 12486
rect 23156 12484 23212 12486
rect 23236 12484 23292 12486
rect 23656 19610 23712 19612
rect 23736 19610 23792 19612
rect 23816 19610 23872 19612
rect 23896 19610 23952 19612
rect 23976 19610 24032 19612
rect 23656 19558 23658 19610
rect 23658 19558 23710 19610
rect 23710 19558 23712 19610
rect 23736 19558 23774 19610
rect 23774 19558 23786 19610
rect 23786 19558 23792 19610
rect 23816 19558 23838 19610
rect 23838 19558 23850 19610
rect 23850 19558 23872 19610
rect 23896 19558 23902 19610
rect 23902 19558 23914 19610
rect 23914 19558 23952 19610
rect 23976 19558 23978 19610
rect 23978 19558 24030 19610
rect 24030 19558 24032 19610
rect 23656 19556 23712 19558
rect 23736 19556 23792 19558
rect 23816 19556 23872 19558
rect 23896 19556 23952 19558
rect 23976 19556 24032 19558
rect 23656 18522 23712 18524
rect 23736 18522 23792 18524
rect 23816 18522 23872 18524
rect 23896 18522 23952 18524
rect 23976 18522 24032 18524
rect 23656 18470 23658 18522
rect 23658 18470 23710 18522
rect 23710 18470 23712 18522
rect 23736 18470 23774 18522
rect 23774 18470 23786 18522
rect 23786 18470 23792 18522
rect 23816 18470 23838 18522
rect 23838 18470 23850 18522
rect 23850 18470 23872 18522
rect 23896 18470 23902 18522
rect 23902 18470 23914 18522
rect 23914 18470 23952 18522
rect 23976 18470 23978 18522
rect 23978 18470 24030 18522
rect 24030 18470 24032 18522
rect 23656 18468 23712 18470
rect 23736 18468 23792 18470
rect 23816 18468 23872 18470
rect 23896 18468 23952 18470
rect 23976 18468 24032 18470
rect 23656 17434 23712 17436
rect 23736 17434 23792 17436
rect 23816 17434 23872 17436
rect 23896 17434 23952 17436
rect 23976 17434 24032 17436
rect 23656 17382 23658 17434
rect 23658 17382 23710 17434
rect 23710 17382 23712 17434
rect 23736 17382 23774 17434
rect 23774 17382 23786 17434
rect 23786 17382 23792 17434
rect 23816 17382 23838 17434
rect 23838 17382 23850 17434
rect 23850 17382 23872 17434
rect 23896 17382 23902 17434
rect 23902 17382 23914 17434
rect 23914 17382 23952 17434
rect 23976 17382 23978 17434
rect 23978 17382 24030 17434
rect 24030 17382 24032 17434
rect 23656 17380 23712 17382
rect 23736 17380 23792 17382
rect 23816 17380 23872 17382
rect 23896 17380 23952 17382
rect 23976 17380 24032 17382
rect 23656 16346 23712 16348
rect 23736 16346 23792 16348
rect 23816 16346 23872 16348
rect 23896 16346 23952 16348
rect 23976 16346 24032 16348
rect 23656 16294 23658 16346
rect 23658 16294 23710 16346
rect 23710 16294 23712 16346
rect 23736 16294 23774 16346
rect 23774 16294 23786 16346
rect 23786 16294 23792 16346
rect 23816 16294 23838 16346
rect 23838 16294 23850 16346
rect 23850 16294 23872 16346
rect 23896 16294 23902 16346
rect 23902 16294 23914 16346
rect 23914 16294 23952 16346
rect 23976 16294 23978 16346
rect 23978 16294 24030 16346
rect 24030 16294 24032 16346
rect 23656 16292 23712 16294
rect 23736 16292 23792 16294
rect 23816 16292 23872 16294
rect 23896 16292 23952 16294
rect 23976 16292 24032 16294
rect 23656 15258 23712 15260
rect 23736 15258 23792 15260
rect 23816 15258 23872 15260
rect 23896 15258 23952 15260
rect 23976 15258 24032 15260
rect 23656 15206 23658 15258
rect 23658 15206 23710 15258
rect 23710 15206 23712 15258
rect 23736 15206 23774 15258
rect 23774 15206 23786 15258
rect 23786 15206 23792 15258
rect 23816 15206 23838 15258
rect 23838 15206 23850 15258
rect 23850 15206 23872 15258
rect 23896 15206 23902 15258
rect 23902 15206 23914 15258
rect 23914 15206 23952 15258
rect 23976 15206 23978 15258
rect 23978 15206 24030 15258
rect 24030 15206 24032 15258
rect 23656 15204 23712 15206
rect 23736 15204 23792 15206
rect 23816 15204 23872 15206
rect 23896 15204 23952 15206
rect 23976 15204 24032 15206
rect 26514 22500 26570 22536
rect 26514 22480 26516 22500
rect 26516 22480 26568 22500
rect 26568 22480 26570 22500
rect 23656 14170 23712 14172
rect 23736 14170 23792 14172
rect 23816 14170 23872 14172
rect 23896 14170 23952 14172
rect 23976 14170 24032 14172
rect 23656 14118 23658 14170
rect 23658 14118 23710 14170
rect 23710 14118 23712 14170
rect 23736 14118 23774 14170
rect 23774 14118 23786 14170
rect 23786 14118 23792 14170
rect 23816 14118 23838 14170
rect 23838 14118 23850 14170
rect 23850 14118 23872 14170
rect 23896 14118 23902 14170
rect 23902 14118 23914 14170
rect 23914 14118 23952 14170
rect 23976 14118 23978 14170
rect 23978 14118 24030 14170
rect 24030 14118 24032 14170
rect 23656 14116 23712 14118
rect 23736 14116 23792 14118
rect 23816 14116 23872 14118
rect 23896 14116 23952 14118
rect 23976 14116 24032 14118
rect 20718 8472 20774 8528
rect 19656 5466 19712 5468
rect 19736 5466 19792 5468
rect 19816 5466 19872 5468
rect 19896 5466 19952 5468
rect 19976 5466 20032 5468
rect 19656 5414 19658 5466
rect 19658 5414 19710 5466
rect 19710 5414 19712 5466
rect 19736 5414 19774 5466
rect 19774 5414 19786 5466
rect 19786 5414 19792 5466
rect 19816 5414 19838 5466
rect 19838 5414 19850 5466
rect 19850 5414 19872 5466
rect 19896 5414 19902 5466
rect 19902 5414 19914 5466
rect 19914 5414 19952 5466
rect 19976 5414 19978 5466
rect 19978 5414 20030 5466
rect 20030 5414 20032 5466
rect 19656 5412 19712 5414
rect 19736 5412 19792 5414
rect 19816 5412 19872 5414
rect 19896 5412 19952 5414
rect 19976 5412 20032 5414
rect 19656 4378 19712 4380
rect 19736 4378 19792 4380
rect 19816 4378 19872 4380
rect 19896 4378 19952 4380
rect 19976 4378 20032 4380
rect 19656 4326 19658 4378
rect 19658 4326 19710 4378
rect 19710 4326 19712 4378
rect 19736 4326 19774 4378
rect 19774 4326 19786 4378
rect 19786 4326 19792 4378
rect 19816 4326 19838 4378
rect 19838 4326 19850 4378
rect 19850 4326 19872 4378
rect 19896 4326 19902 4378
rect 19902 4326 19914 4378
rect 19914 4326 19952 4378
rect 19976 4326 19978 4378
rect 19978 4326 20030 4378
rect 20030 4326 20032 4378
rect 19656 4324 19712 4326
rect 19736 4324 19792 4326
rect 19816 4324 19872 4326
rect 19896 4324 19952 4326
rect 19976 4324 20032 4326
rect 20994 6704 21050 6760
rect 20902 6296 20958 6352
rect 22916 11450 22972 11452
rect 22996 11450 23052 11452
rect 23076 11450 23132 11452
rect 23156 11450 23212 11452
rect 23236 11450 23292 11452
rect 22916 11398 22918 11450
rect 22918 11398 22970 11450
rect 22970 11398 22972 11450
rect 22996 11398 23034 11450
rect 23034 11398 23046 11450
rect 23046 11398 23052 11450
rect 23076 11398 23098 11450
rect 23098 11398 23110 11450
rect 23110 11398 23132 11450
rect 23156 11398 23162 11450
rect 23162 11398 23174 11450
rect 23174 11398 23212 11450
rect 23236 11398 23238 11450
rect 23238 11398 23290 11450
rect 23290 11398 23292 11450
rect 22916 11396 22972 11398
rect 22996 11396 23052 11398
rect 23076 11396 23132 11398
rect 23156 11396 23212 11398
rect 23236 11396 23292 11398
rect 22916 10362 22972 10364
rect 22996 10362 23052 10364
rect 23076 10362 23132 10364
rect 23156 10362 23212 10364
rect 23236 10362 23292 10364
rect 22916 10310 22918 10362
rect 22918 10310 22970 10362
rect 22970 10310 22972 10362
rect 22996 10310 23034 10362
rect 23034 10310 23046 10362
rect 23046 10310 23052 10362
rect 23076 10310 23098 10362
rect 23098 10310 23110 10362
rect 23110 10310 23132 10362
rect 23156 10310 23162 10362
rect 23162 10310 23174 10362
rect 23174 10310 23212 10362
rect 23236 10310 23238 10362
rect 23238 10310 23290 10362
rect 23290 10310 23292 10362
rect 22916 10308 22972 10310
rect 22996 10308 23052 10310
rect 23076 10308 23132 10310
rect 23156 10308 23212 10310
rect 23236 10308 23292 10310
rect 21638 7268 21694 7304
rect 21638 7248 21640 7268
rect 21640 7248 21692 7268
rect 21692 7248 21694 7268
rect 22098 6316 22154 6352
rect 22098 6296 22100 6316
rect 22100 6296 22152 6316
rect 22152 6296 22154 6316
rect 22916 9274 22972 9276
rect 22996 9274 23052 9276
rect 23076 9274 23132 9276
rect 23156 9274 23212 9276
rect 23236 9274 23292 9276
rect 22916 9222 22918 9274
rect 22918 9222 22970 9274
rect 22970 9222 22972 9274
rect 22996 9222 23034 9274
rect 23034 9222 23046 9274
rect 23046 9222 23052 9274
rect 23076 9222 23098 9274
rect 23098 9222 23110 9274
rect 23110 9222 23132 9274
rect 23156 9222 23162 9274
rect 23162 9222 23174 9274
rect 23174 9222 23212 9274
rect 23236 9222 23238 9274
rect 23238 9222 23290 9274
rect 23290 9222 23292 9274
rect 22916 9220 22972 9222
rect 22996 9220 23052 9222
rect 23076 9220 23132 9222
rect 23156 9220 23212 9222
rect 23236 9220 23292 9222
rect 23656 13082 23712 13084
rect 23736 13082 23792 13084
rect 23816 13082 23872 13084
rect 23896 13082 23952 13084
rect 23976 13082 24032 13084
rect 23656 13030 23658 13082
rect 23658 13030 23710 13082
rect 23710 13030 23712 13082
rect 23736 13030 23774 13082
rect 23774 13030 23786 13082
rect 23786 13030 23792 13082
rect 23816 13030 23838 13082
rect 23838 13030 23850 13082
rect 23850 13030 23872 13082
rect 23896 13030 23902 13082
rect 23902 13030 23914 13082
rect 23914 13030 23952 13082
rect 23976 13030 23978 13082
rect 23978 13030 24030 13082
rect 24030 13030 24032 13082
rect 23656 13028 23712 13030
rect 23736 13028 23792 13030
rect 23816 13028 23872 13030
rect 23896 13028 23952 13030
rect 23976 13028 24032 13030
rect 23656 11994 23712 11996
rect 23736 11994 23792 11996
rect 23816 11994 23872 11996
rect 23896 11994 23952 11996
rect 23976 11994 24032 11996
rect 23656 11942 23658 11994
rect 23658 11942 23710 11994
rect 23710 11942 23712 11994
rect 23736 11942 23774 11994
rect 23774 11942 23786 11994
rect 23786 11942 23792 11994
rect 23816 11942 23838 11994
rect 23838 11942 23850 11994
rect 23850 11942 23872 11994
rect 23896 11942 23902 11994
rect 23902 11942 23914 11994
rect 23914 11942 23952 11994
rect 23976 11942 23978 11994
rect 23978 11942 24030 11994
rect 24030 11942 24032 11994
rect 23656 11940 23712 11942
rect 23736 11940 23792 11942
rect 23816 11940 23872 11942
rect 23896 11940 23952 11942
rect 23976 11940 24032 11942
rect 23656 10906 23712 10908
rect 23736 10906 23792 10908
rect 23816 10906 23872 10908
rect 23896 10906 23952 10908
rect 23976 10906 24032 10908
rect 23656 10854 23658 10906
rect 23658 10854 23710 10906
rect 23710 10854 23712 10906
rect 23736 10854 23774 10906
rect 23774 10854 23786 10906
rect 23786 10854 23792 10906
rect 23816 10854 23838 10906
rect 23838 10854 23850 10906
rect 23850 10854 23872 10906
rect 23896 10854 23902 10906
rect 23902 10854 23914 10906
rect 23914 10854 23952 10906
rect 23976 10854 23978 10906
rect 23978 10854 24030 10906
rect 24030 10854 24032 10906
rect 23656 10852 23712 10854
rect 23736 10852 23792 10854
rect 23816 10852 23872 10854
rect 23896 10852 23952 10854
rect 23976 10852 24032 10854
rect 23656 9818 23712 9820
rect 23736 9818 23792 9820
rect 23816 9818 23872 9820
rect 23896 9818 23952 9820
rect 23976 9818 24032 9820
rect 23656 9766 23658 9818
rect 23658 9766 23710 9818
rect 23710 9766 23712 9818
rect 23736 9766 23774 9818
rect 23774 9766 23786 9818
rect 23786 9766 23792 9818
rect 23816 9766 23838 9818
rect 23838 9766 23850 9818
rect 23850 9766 23872 9818
rect 23896 9766 23902 9818
rect 23902 9766 23914 9818
rect 23914 9766 23952 9818
rect 23976 9766 23978 9818
rect 23978 9766 24030 9818
rect 24030 9766 24032 9818
rect 23656 9764 23712 9766
rect 23736 9764 23792 9766
rect 23816 9764 23872 9766
rect 23896 9764 23952 9766
rect 23976 9764 24032 9766
rect 25962 13640 26018 13696
rect 22916 8186 22972 8188
rect 22996 8186 23052 8188
rect 23076 8186 23132 8188
rect 23156 8186 23212 8188
rect 23236 8186 23292 8188
rect 22916 8134 22918 8186
rect 22918 8134 22970 8186
rect 22970 8134 22972 8186
rect 22996 8134 23034 8186
rect 23034 8134 23046 8186
rect 23046 8134 23052 8186
rect 23076 8134 23098 8186
rect 23098 8134 23110 8186
rect 23110 8134 23132 8186
rect 23156 8134 23162 8186
rect 23162 8134 23174 8186
rect 23174 8134 23212 8186
rect 23236 8134 23238 8186
rect 23238 8134 23290 8186
rect 23290 8134 23292 8186
rect 22916 8132 22972 8134
rect 22996 8132 23052 8134
rect 23076 8132 23132 8134
rect 23156 8132 23212 8134
rect 23236 8132 23292 8134
rect 22916 7098 22972 7100
rect 22996 7098 23052 7100
rect 23076 7098 23132 7100
rect 23156 7098 23212 7100
rect 23236 7098 23292 7100
rect 22916 7046 22918 7098
rect 22918 7046 22970 7098
rect 22970 7046 22972 7098
rect 22996 7046 23034 7098
rect 23034 7046 23046 7098
rect 23046 7046 23052 7098
rect 23076 7046 23098 7098
rect 23098 7046 23110 7098
rect 23110 7046 23132 7098
rect 23156 7046 23162 7098
rect 23162 7046 23174 7098
rect 23174 7046 23212 7098
rect 23236 7046 23238 7098
rect 23238 7046 23290 7098
rect 23290 7046 23292 7098
rect 22916 7044 22972 7046
rect 22996 7044 23052 7046
rect 23076 7044 23132 7046
rect 23156 7044 23212 7046
rect 23236 7044 23292 7046
rect 19656 3290 19712 3292
rect 19736 3290 19792 3292
rect 19816 3290 19872 3292
rect 19896 3290 19952 3292
rect 19976 3290 20032 3292
rect 19656 3238 19658 3290
rect 19658 3238 19710 3290
rect 19710 3238 19712 3290
rect 19736 3238 19774 3290
rect 19774 3238 19786 3290
rect 19786 3238 19792 3290
rect 19816 3238 19838 3290
rect 19838 3238 19850 3290
rect 19850 3238 19872 3290
rect 19896 3238 19902 3290
rect 19902 3238 19914 3290
rect 19914 3238 19952 3290
rect 19976 3238 19978 3290
rect 19978 3238 20030 3290
rect 20030 3238 20032 3290
rect 19656 3236 19712 3238
rect 19736 3236 19792 3238
rect 19816 3236 19872 3238
rect 19896 3236 19952 3238
rect 19976 3236 20032 3238
rect 23656 8730 23712 8732
rect 23736 8730 23792 8732
rect 23816 8730 23872 8732
rect 23896 8730 23952 8732
rect 23976 8730 24032 8732
rect 23656 8678 23658 8730
rect 23658 8678 23710 8730
rect 23710 8678 23712 8730
rect 23736 8678 23774 8730
rect 23774 8678 23786 8730
rect 23786 8678 23792 8730
rect 23816 8678 23838 8730
rect 23838 8678 23850 8730
rect 23850 8678 23872 8730
rect 23896 8678 23902 8730
rect 23902 8678 23914 8730
rect 23914 8678 23952 8730
rect 23976 8678 23978 8730
rect 23978 8678 24030 8730
rect 24030 8678 24032 8730
rect 23656 8676 23712 8678
rect 23736 8676 23792 8678
rect 23816 8676 23872 8678
rect 23896 8676 23952 8678
rect 23976 8676 24032 8678
rect 23656 7642 23712 7644
rect 23736 7642 23792 7644
rect 23816 7642 23872 7644
rect 23896 7642 23952 7644
rect 23976 7642 24032 7644
rect 23656 7590 23658 7642
rect 23658 7590 23710 7642
rect 23710 7590 23712 7642
rect 23736 7590 23774 7642
rect 23774 7590 23786 7642
rect 23786 7590 23792 7642
rect 23816 7590 23838 7642
rect 23838 7590 23850 7642
rect 23850 7590 23872 7642
rect 23896 7590 23902 7642
rect 23902 7590 23914 7642
rect 23914 7590 23952 7642
rect 23976 7590 23978 7642
rect 23978 7590 24030 7642
rect 24030 7590 24032 7642
rect 23656 7588 23712 7590
rect 23736 7588 23792 7590
rect 23816 7588 23872 7590
rect 23896 7588 23952 7590
rect 23976 7588 24032 7590
rect 23656 6554 23712 6556
rect 23736 6554 23792 6556
rect 23816 6554 23872 6556
rect 23896 6554 23952 6556
rect 23976 6554 24032 6556
rect 23656 6502 23658 6554
rect 23658 6502 23710 6554
rect 23710 6502 23712 6554
rect 23736 6502 23774 6554
rect 23774 6502 23786 6554
rect 23786 6502 23792 6554
rect 23816 6502 23838 6554
rect 23838 6502 23850 6554
rect 23850 6502 23872 6554
rect 23896 6502 23902 6554
rect 23902 6502 23914 6554
rect 23914 6502 23952 6554
rect 23976 6502 23978 6554
rect 23978 6502 24030 6554
rect 24030 6502 24032 6554
rect 23656 6500 23712 6502
rect 23736 6500 23792 6502
rect 23816 6500 23872 6502
rect 23896 6500 23952 6502
rect 23976 6500 24032 6502
rect 22916 6010 22972 6012
rect 22996 6010 23052 6012
rect 23076 6010 23132 6012
rect 23156 6010 23212 6012
rect 23236 6010 23292 6012
rect 22916 5958 22918 6010
rect 22918 5958 22970 6010
rect 22970 5958 22972 6010
rect 22996 5958 23034 6010
rect 23034 5958 23046 6010
rect 23046 5958 23052 6010
rect 23076 5958 23098 6010
rect 23098 5958 23110 6010
rect 23110 5958 23132 6010
rect 23156 5958 23162 6010
rect 23162 5958 23174 6010
rect 23174 5958 23212 6010
rect 23236 5958 23238 6010
rect 23238 5958 23290 6010
rect 23290 5958 23292 6010
rect 22916 5956 22972 5958
rect 22996 5956 23052 5958
rect 23076 5956 23132 5958
rect 23156 5956 23212 5958
rect 23236 5956 23292 5958
rect 23656 5466 23712 5468
rect 23736 5466 23792 5468
rect 23816 5466 23872 5468
rect 23896 5466 23952 5468
rect 23976 5466 24032 5468
rect 23656 5414 23658 5466
rect 23658 5414 23710 5466
rect 23710 5414 23712 5466
rect 23736 5414 23774 5466
rect 23774 5414 23786 5466
rect 23786 5414 23792 5466
rect 23816 5414 23838 5466
rect 23838 5414 23850 5466
rect 23850 5414 23872 5466
rect 23896 5414 23902 5466
rect 23902 5414 23914 5466
rect 23914 5414 23952 5466
rect 23976 5414 23978 5466
rect 23978 5414 24030 5466
rect 24030 5414 24032 5466
rect 23656 5412 23712 5414
rect 23736 5412 23792 5414
rect 23816 5412 23872 5414
rect 23896 5412 23952 5414
rect 23976 5412 24032 5414
rect 22916 4922 22972 4924
rect 22996 4922 23052 4924
rect 23076 4922 23132 4924
rect 23156 4922 23212 4924
rect 23236 4922 23292 4924
rect 22916 4870 22918 4922
rect 22918 4870 22970 4922
rect 22970 4870 22972 4922
rect 22996 4870 23034 4922
rect 23034 4870 23046 4922
rect 23046 4870 23052 4922
rect 23076 4870 23098 4922
rect 23098 4870 23110 4922
rect 23110 4870 23132 4922
rect 23156 4870 23162 4922
rect 23162 4870 23174 4922
rect 23174 4870 23212 4922
rect 23236 4870 23238 4922
rect 23238 4870 23290 4922
rect 23290 4870 23292 4922
rect 22916 4868 22972 4870
rect 22996 4868 23052 4870
rect 23076 4868 23132 4870
rect 23156 4868 23212 4870
rect 23236 4868 23292 4870
rect 26146 9560 26202 9616
rect 25410 6296 25466 6352
rect 26514 7540 26570 7576
rect 26514 7520 26516 7540
rect 26516 7520 26568 7540
rect 26568 7520 26570 7540
rect 26330 7248 26386 7304
rect 25962 6316 26018 6352
rect 25962 6296 25964 6316
rect 25964 6296 26016 6316
rect 26016 6296 26018 6316
rect 22916 3834 22972 3836
rect 22996 3834 23052 3836
rect 23076 3834 23132 3836
rect 23156 3834 23212 3836
rect 23236 3834 23292 3836
rect 22916 3782 22918 3834
rect 22918 3782 22970 3834
rect 22970 3782 22972 3834
rect 22996 3782 23034 3834
rect 23034 3782 23046 3834
rect 23046 3782 23052 3834
rect 23076 3782 23098 3834
rect 23098 3782 23110 3834
rect 23110 3782 23132 3834
rect 23156 3782 23162 3834
rect 23162 3782 23174 3834
rect 23174 3782 23212 3834
rect 23236 3782 23238 3834
rect 23238 3782 23290 3834
rect 23290 3782 23292 3834
rect 22916 3780 22972 3782
rect 22996 3780 23052 3782
rect 23076 3780 23132 3782
rect 23156 3780 23212 3782
rect 23236 3780 23292 3782
rect 23656 4378 23712 4380
rect 23736 4378 23792 4380
rect 23816 4378 23872 4380
rect 23896 4378 23952 4380
rect 23976 4378 24032 4380
rect 23656 4326 23658 4378
rect 23658 4326 23710 4378
rect 23710 4326 23712 4378
rect 23736 4326 23774 4378
rect 23774 4326 23786 4378
rect 23786 4326 23792 4378
rect 23816 4326 23838 4378
rect 23838 4326 23850 4378
rect 23850 4326 23872 4378
rect 23896 4326 23902 4378
rect 23902 4326 23914 4378
rect 23914 4326 23952 4378
rect 23976 4326 23978 4378
rect 23978 4326 24030 4378
rect 24030 4326 24032 4378
rect 23656 4324 23712 4326
rect 23736 4324 23792 4326
rect 23816 4324 23872 4326
rect 23896 4324 23952 4326
rect 23976 4324 24032 4326
rect 23656 3290 23712 3292
rect 23736 3290 23792 3292
rect 23816 3290 23872 3292
rect 23896 3290 23952 3292
rect 23976 3290 24032 3292
rect 23656 3238 23658 3290
rect 23658 3238 23710 3290
rect 23710 3238 23712 3290
rect 23736 3238 23774 3290
rect 23774 3238 23786 3290
rect 23786 3238 23792 3290
rect 23816 3238 23838 3290
rect 23838 3238 23850 3290
rect 23850 3238 23872 3290
rect 23896 3238 23902 3290
rect 23902 3238 23914 3290
rect 23914 3238 23952 3290
rect 23976 3238 23978 3290
rect 23978 3238 24030 3290
rect 24030 3238 24032 3290
rect 23656 3236 23712 3238
rect 23736 3236 23792 3238
rect 23816 3236 23872 3238
rect 23896 3236 23952 3238
rect 23976 3236 24032 3238
rect 22916 2746 22972 2748
rect 22996 2746 23052 2748
rect 23076 2746 23132 2748
rect 23156 2746 23212 2748
rect 23236 2746 23292 2748
rect 22916 2694 22918 2746
rect 22918 2694 22970 2746
rect 22970 2694 22972 2746
rect 22996 2694 23034 2746
rect 23034 2694 23046 2746
rect 23046 2694 23052 2746
rect 23076 2694 23098 2746
rect 23098 2694 23110 2746
rect 23110 2694 23132 2746
rect 23156 2694 23162 2746
rect 23162 2694 23174 2746
rect 23174 2694 23212 2746
rect 23236 2694 23238 2746
rect 23238 2694 23290 2746
rect 23290 2694 23292 2746
rect 22916 2692 22972 2694
rect 22996 2692 23052 2694
rect 23076 2692 23132 2694
rect 23156 2692 23212 2694
rect 23236 2692 23292 2694
rect 19656 2202 19712 2204
rect 19736 2202 19792 2204
rect 19816 2202 19872 2204
rect 19896 2202 19952 2204
rect 19976 2202 20032 2204
rect 19656 2150 19658 2202
rect 19658 2150 19710 2202
rect 19710 2150 19712 2202
rect 19736 2150 19774 2202
rect 19774 2150 19786 2202
rect 19786 2150 19792 2202
rect 19816 2150 19838 2202
rect 19838 2150 19850 2202
rect 19850 2150 19872 2202
rect 19896 2150 19902 2202
rect 19902 2150 19914 2202
rect 19914 2150 19952 2202
rect 19976 2150 19978 2202
rect 19978 2150 20030 2202
rect 20030 2150 20032 2202
rect 19656 2148 19712 2150
rect 19736 2148 19792 2150
rect 19816 2148 19872 2150
rect 19896 2148 19952 2150
rect 19976 2148 20032 2150
rect 23656 2202 23712 2204
rect 23736 2202 23792 2204
rect 23816 2202 23872 2204
rect 23896 2202 23952 2204
rect 23976 2202 24032 2204
rect 23656 2150 23658 2202
rect 23658 2150 23710 2202
rect 23710 2150 23712 2202
rect 23736 2150 23774 2202
rect 23774 2150 23786 2202
rect 23786 2150 23792 2202
rect 23816 2150 23838 2202
rect 23838 2150 23850 2202
rect 23850 2150 23872 2202
rect 23896 2150 23902 2202
rect 23902 2150 23914 2202
rect 23914 2150 23952 2202
rect 23976 2150 23978 2202
rect 23978 2150 24030 2202
rect 24030 2150 24032 2202
rect 23656 2148 23712 2150
rect 23736 2148 23792 2150
rect 23816 2148 23872 2150
rect 23896 2148 23952 2150
rect 23976 2148 24032 2150
<< metal3 >>
rect 2906 27776 3302 27777
rect 2906 27712 2912 27776
rect 2976 27712 2992 27776
rect 3056 27712 3072 27776
rect 3136 27712 3152 27776
rect 3216 27712 3232 27776
rect 3296 27712 3302 27776
rect 2906 27711 3302 27712
rect 6906 27776 7302 27777
rect 6906 27712 6912 27776
rect 6976 27712 6992 27776
rect 7056 27712 7072 27776
rect 7136 27712 7152 27776
rect 7216 27712 7232 27776
rect 7296 27712 7302 27776
rect 6906 27711 7302 27712
rect 10906 27776 11302 27777
rect 10906 27712 10912 27776
rect 10976 27712 10992 27776
rect 11056 27712 11072 27776
rect 11136 27712 11152 27776
rect 11216 27712 11232 27776
rect 11296 27712 11302 27776
rect 10906 27711 11302 27712
rect 14906 27776 15302 27777
rect 14906 27712 14912 27776
rect 14976 27712 14992 27776
rect 15056 27712 15072 27776
rect 15136 27712 15152 27776
rect 15216 27712 15232 27776
rect 15296 27712 15302 27776
rect 14906 27711 15302 27712
rect 18906 27776 19302 27777
rect 18906 27712 18912 27776
rect 18976 27712 18992 27776
rect 19056 27712 19072 27776
rect 19136 27712 19152 27776
rect 19216 27712 19232 27776
rect 19296 27712 19302 27776
rect 18906 27711 19302 27712
rect 22906 27776 23302 27777
rect 22906 27712 22912 27776
rect 22976 27712 22992 27776
rect 23056 27712 23072 27776
rect 23136 27712 23152 27776
rect 23216 27712 23232 27776
rect 23296 27712 23302 27776
rect 22906 27711 23302 27712
rect 3646 27232 4042 27233
rect 3646 27168 3652 27232
rect 3716 27168 3732 27232
rect 3796 27168 3812 27232
rect 3876 27168 3892 27232
rect 3956 27168 3972 27232
rect 4036 27168 4042 27232
rect 3646 27167 4042 27168
rect 7646 27232 8042 27233
rect 7646 27168 7652 27232
rect 7716 27168 7732 27232
rect 7796 27168 7812 27232
rect 7876 27168 7892 27232
rect 7956 27168 7972 27232
rect 8036 27168 8042 27232
rect 7646 27167 8042 27168
rect 11646 27232 12042 27233
rect 11646 27168 11652 27232
rect 11716 27168 11732 27232
rect 11796 27168 11812 27232
rect 11876 27168 11892 27232
rect 11956 27168 11972 27232
rect 12036 27168 12042 27232
rect 11646 27167 12042 27168
rect 15646 27232 16042 27233
rect 15646 27168 15652 27232
rect 15716 27168 15732 27232
rect 15796 27168 15812 27232
rect 15876 27168 15892 27232
rect 15956 27168 15972 27232
rect 16036 27168 16042 27232
rect 15646 27167 16042 27168
rect 19646 27232 20042 27233
rect 19646 27168 19652 27232
rect 19716 27168 19732 27232
rect 19796 27168 19812 27232
rect 19876 27168 19892 27232
rect 19956 27168 19972 27232
rect 20036 27168 20042 27232
rect 19646 27167 20042 27168
rect 23646 27232 24042 27233
rect 23646 27168 23652 27232
rect 23716 27168 23732 27232
rect 23796 27168 23812 27232
rect 23876 27168 23892 27232
rect 23956 27168 23972 27232
rect 24036 27168 24042 27232
rect 23646 27167 24042 27168
rect 10174 26828 10180 26892
rect 10244 26890 10250 26892
rect 10869 26890 10935 26893
rect 10244 26888 10935 26890
rect 10244 26832 10874 26888
rect 10930 26832 10935 26888
rect 10244 26830 10935 26832
rect 10244 26828 10250 26830
rect 10869 26827 10935 26830
rect 2906 26688 3302 26689
rect 0 26618 800 26648
rect 2906 26624 2912 26688
rect 2976 26624 2992 26688
rect 3056 26624 3072 26688
rect 3136 26624 3152 26688
rect 3216 26624 3232 26688
rect 3296 26624 3302 26688
rect 2906 26623 3302 26624
rect 6906 26688 7302 26689
rect 6906 26624 6912 26688
rect 6976 26624 6992 26688
rect 7056 26624 7072 26688
rect 7136 26624 7152 26688
rect 7216 26624 7232 26688
rect 7296 26624 7302 26688
rect 6906 26623 7302 26624
rect 10906 26688 11302 26689
rect 10906 26624 10912 26688
rect 10976 26624 10992 26688
rect 11056 26624 11072 26688
rect 11136 26624 11152 26688
rect 11216 26624 11232 26688
rect 11296 26624 11302 26688
rect 10906 26623 11302 26624
rect 14906 26688 15302 26689
rect 14906 26624 14912 26688
rect 14976 26624 14992 26688
rect 15056 26624 15072 26688
rect 15136 26624 15152 26688
rect 15216 26624 15232 26688
rect 15296 26624 15302 26688
rect 14906 26623 15302 26624
rect 18906 26688 19302 26689
rect 18906 26624 18912 26688
rect 18976 26624 18992 26688
rect 19056 26624 19072 26688
rect 19136 26624 19152 26688
rect 19216 26624 19232 26688
rect 19296 26624 19302 26688
rect 18906 26623 19302 26624
rect 22906 26688 23302 26689
rect 22906 26624 22912 26688
rect 22976 26624 22992 26688
rect 23056 26624 23072 26688
rect 23136 26624 23152 26688
rect 23216 26624 23232 26688
rect 23296 26624 23302 26688
rect 22906 26623 23302 26624
rect 0 26558 1778 26618
rect 0 26528 800 26558
rect 1718 26482 1778 26558
rect 3417 26482 3483 26485
rect 1718 26480 3483 26482
rect 1718 26424 3422 26480
rect 3478 26424 3483 26480
rect 1718 26422 3483 26424
rect 3417 26419 3483 26422
rect 3646 26144 4042 26145
rect 3646 26080 3652 26144
rect 3716 26080 3732 26144
rect 3796 26080 3812 26144
rect 3876 26080 3892 26144
rect 3956 26080 3972 26144
rect 4036 26080 4042 26144
rect 3646 26079 4042 26080
rect 7646 26144 8042 26145
rect 7646 26080 7652 26144
rect 7716 26080 7732 26144
rect 7796 26080 7812 26144
rect 7876 26080 7892 26144
rect 7956 26080 7972 26144
rect 8036 26080 8042 26144
rect 7646 26079 8042 26080
rect 11646 26144 12042 26145
rect 11646 26080 11652 26144
rect 11716 26080 11732 26144
rect 11796 26080 11812 26144
rect 11876 26080 11892 26144
rect 11956 26080 11972 26144
rect 12036 26080 12042 26144
rect 11646 26079 12042 26080
rect 15646 26144 16042 26145
rect 15646 26080 15652 26144
rect 15716 26080 15732 26144
rect 15796 26080 15812 26144
rect 15876 26080 15892 26144
rect 15956 26080 15972 26144
rect 16036 26080 16042 26144
rect 15646 26079 16042 26080
rect 19646 26144 20042 26145
rect 19646 26080 19652 26144
rect 19716 26080 19732 26144
rect 19796 26080 19812 26144
rect 19876 26080 19892 26144
rect 19956 26080 19972 26144
rect 20036 26080 20042 26144
rect 19646 26079 20042 26080
rect 23646 26144 24042 26145
rect 23646 26080 23652 26144
rect 23716 26080 23732 26144
rect 23796 26080 23812 26144
rect 23876 26080 23892 26144
rect 23956 26080 23972 26144
rect 24036 26080 24042 26144
rect 23646 26079 24042 26080
rect 2906 25600 3302 25601
rect 2906 25536 2912 25600
rect 2976 25536 2992 25600
rect 3056 25536 3072 25600
rect 3136 25536 3152 25600
rect 3216 25536 3232 25600
rect 3296 25536 3302 25600
rect 2906 25535 3302 25536
rect 6906 25600 7302 25601
rect 6906 25536 6912 25600
rect 6976 25536 6992 25600
rect 7056 25536 7072 25600
rect 7136 25536 7152 25600
rect 7216 25536 7232 25600
rect 7296 25536 7302 25600
rect 6906 25535 7302 25536
rect 10906 25600 11302 25601
rect 10906 25536 10912 25600
rect 10976 25536 10992 25600
rect 11056 25536 11072 25600
rect 11136 25536 11152 25600
rect 11216 25536 11232 25600
rect 11296 25536 11302 25600
rect 10906 25535 11302 25536
rect 14906 25600 15302 25601
rect 14906 25536 14912 25600
rect 14976 25536 14992 25600
rect 15056 25536 15072 25600
rect 15136 25536 15152 25600
rect 15216 25536 15232 25600
rect 15296 25536 15302 25600
rect 14906 25535 15302 25536
rect 18906 25600 19302 25601
rect 18906 25536 18912 25600
rect 18976 25536 18992 25600
rect 19056 25536 19072 25600
rect 19136 25536 19152 25600
rect 19216 25536 19232 25600
rect 19296 25536 19302 25600
rect 18906 25535 19302 25536
rect 22906 25600 23302 25601
rect 22906 25536 22912 25600
rect 22976 25536 22992 25600
rect 23056 25536 23072 25600
rect 23136 25536 23152 25600
rect 23216 25536 23232 25600
rect 23296 25536 23302 25600
rect 22906 25535 23302 25536
rect 3646 25056 4042 25057
rect 3646 24992 3652 25056
rect 3716 24992 3732 25056
rect 3796 24992 3812 25056
rect 3876 24992 3892 25056
rect 3956 24992 3972 25056
rect 4036 24992 4042 25056
rect 3646 24991 4042 24992
rect 7646 25056 8042 25057
rect 7646 24992 7652 25056
rect 7716 24992 7732 25056
rect 7796 24992 7812 25056
rect 7876 24992 7892 25056
rect 7956 24992 7972 25056
rect 8036 24992 8042 25056
rect 7646 24991 8042 24992
rect 11646 25056 12042 25057
rect 11646 24992 11652 25056
rect 11716 24992 11732 25056
rect 11796 24992 11812 25056
rect 11876 24992 11892 25056
rect 11956 24992 11972 25056
rect 12036 24992 12042 25056
rect 11646 24991 12042 24992
rect 15646 25056 16042 25057
rect 15646 24992 15652 25056
rect 15716 24992 15732 25056
rect 15796 24992 15812 25056
rect 15876 24992 15892 25056
rect 15956 24992 15972 25056
rect 16036 24992 16042 25056
rect 15646 24991 16042 24992
rect 19646 25056 20042 25057
rect 19646 24992 19652 25056
rect 19716 24992 19732 25056
rect 19796 24992 19812 25056
rect 19876 24992 19892 25056
rect 19956 24992 19972 25056
rect 20036 24992 20042 25056
rect 19646 24991 20042 24992
rect 23646 25056 24042 25057
rect 23646 24992 23652 25056
rect 23716 24992 23732 25056
rect 23796 24992 23812 25056
rect 23876 24992 23892 25056
rect 23956 24992 23972 25056
rect 24036 24992 24042 25056
rect 23646 24991 24042 24992
rect 17534 24924 17540 24988
rect 17604 24986 17610 24988
rect 17677 24986 17743 24989
rect 17604 24984 17743 24986
rect 17604 24928 17682 24984
rect 17738 24928 17743 24984
rect 17604 24926 17743 24928
rect 17604 24924 17610 24926
rect 17677 24923 17743 24926
rect 24342 24924 24348 24988
rect 24412 24986 24418 24988
rect 24485 24986 24551 24989
rect 24412 24984 24551 24986
rect 24412 24928 24490 24984
rect 24546 24928 24551 24984
rect 24412 24926 24551 24928
rect 24412 24924 24418 24926
rect 24485 24923 24551 24926
rect 2906 24512 3302 24513
rect 2906 24448 2912 24512
rect 2976 24448 2992 24512
rect 3056 24448 3072 24512
rect 3136 24448 3152 24512
rect 3216 24448 3232 24512
rect 3296 24448 3302 24512
rect 2906 24447 3302 24448
rect 6906 24512 7302 24513
rect 6906 24448 6912 24512
rect 6976 24448 6992 24512
rect 7056 24448 7072 24512
rect 7136 24448 7152 24512
rect 7216 24448 7232 24512
rect 7296 24448 7302 24512
rect 6906 24447 7302 24448
rect 10906 24512 11302 24513
rect 10906 24448 10912 24512
rect 10976 24448 10992 24512
rect 11056 24448 11072 24512
rect 11136 24448 11152 24512
rect 11216 24448 11232 24512
rect 11296 24448 11302 24512
rect 10906 24447 11302 24448
rect 14906 24512 15302 24513
rect 14906 24448 14912 24512
rect 14976 24448 14992 24512
rect 15056 24448 15072 24512
rect 15136 24448 15152 24512
rect 15216 24448 15232 24512
rect 15296 24448 15302 24512
rect 14906 24447 15302 24448
rect 18906 24512 19302 24513
rect 18906 24448 18912 24512
rect 18976 24448 18992 24512
rect 19056 24448 19072 24512
rect 19136 24448 19152 24512
rect 19216 24448 19232 24512
rect 19296 24448 19302 24512
rect 18906 24447 19302 24448
rect 22906 24512 23302 24513
rect 22906 24448 22912 24512
rect 22976 24448 22992 24512
rect 23056 24448 23072 24512
rect 23136 24448 23152 24512
rect 23216 24448 23232 24512
rect 23296 24448 23302 24512
rect 22906 24447 23302 24448
rect 3646 23968 4042 23969
rect 3646 23904 3652 23968
rect 3716 23904 3732 23968
rect 3796 23904 3812 23968
rect 3876 23904 3892 23968
rect 3956 23904 3972 23968
rect 4036 23904 4042 23968
rect 3646 23903 4042 23904
rect 7646 23968 8042 23969
rect 7646 23904 7652 23968
rect 7716 23904 7732 23968
rect 7796 23904 7812 23968
rect 7876 23904 7892 23968
rect 7956 23904 7972 23968
rect 8036 23904 8042 23968
rect 7646 23903 8042 23904
rect 11646 23968 12042 23969
rect 11646 23904 11652 23968
rect 11716 23904 11732 23968
rect 11796 23904 11812 23968
rect 11876 23904 11892 23968
rect 11956 23904 11972 23968
rect 12036 23904 12042 23968
rect 11646 23903 12042 23904
rect 15646 23968 16042 23969
rect 15646 23904 15652 23968
rect 15716 23904 15732 23968
rect 15796 23904 15812 23968
rect 15876 23904 15892 23968
rect 15956 23904 15972 23968
rect 16036 23904 16042 23968
rect 15646 23903 16042 23904
rect 19646 23968 20042 23969
rect 19646 23904 19652 23968
rect 19716 23904 19732 23968
rect 19796 23904 19812 23968
rect 19876 23904 19892 23968
rect 19956 23904 19972 23968
rect 20036 23904 20042 23968
rect 19646 23903 20042 23904
rect 23646 23968 24042 23969
rect 23646 23904 23652 23968
rect 23716 23904 23732 23968
rect 23796 23904 23812 23968
rect 23876 23904 23892 23968
rect 23956 23904 23972 23968
rect 24036 23904 24042 23968
rect 23646 23903 24042 23904
rect 2906 23424 3302 23425
rect 2906 23360 2912 23424
rect 2976 23360 2992 23424
rect 3056 23360 3072 23424
rect 3136 23360 3152 23424
rect 3216 23360 3232 23424
rect 3296 23360 3302 23424
rect 2906 23359 3302 23360
rect 6906 23424 7302 23425
rect 6906 23360 6912 23424
rect 6976 23360 6992 23424
rect 7056 23360 7072 23424
rect 7136 23360 7152 23424
rect 7216 23360 7232 23424
rect 7296 23360 7302 23424
rect 6906 23359 7302 23360
rect 10906 23424 11302 23425
rect 10906 23360 10912 23424
rect 10976 23360 10992 23424
rect 11056 23360 11072 23424
rect 11136 23360 11152 23424
rect 11216 23360 11232 23424
rect 11296 23360 11302 23424
rect 10906 23359 11302 23360
rect 14906 23424 15302 23425
rect 14906 23360 14912 23424
rect 14976 23360 14992 23424
rect 15056 23360 15072 23424
rect 15136 23360 15152 23424
rect 15216 23360 15232 23424
rect 15296 23360 15302 23424
rect 14906 23359 15302 23360
rect 18906 23424 19302 23425
rect 18906 23360 18912 23424
rect 18976 23360 18992 23424
rect 19056 23360 19072 23424
rect 19136 23360 19152 23424
rect 19216 23360 19232 23424
rect 19296 23360 19302 23424
rect 18906 23359 19302 23360
rect 22906 23424 23302 23425
rect 22906 23360 22912 23424
rect 22976 23360 22992 23424
rect 23056 23360 23072 23424
rect 23136 23360 23152 23424
rect 23216 23360 23232 23424
rect 23296 23360 23302 23424
rect 22906 23359 23302 23360
rect 10869 23082 10935 23085
rect 12893 23082 12959 23085
rect 10869 23080 12959 23082
rect 10869 23024 10874 23080
rect 10930 23024 12898 23080
rect 12954 23024 12959 23080
rect 10869 23022 12959 23024
rect 10869 23019 10935 23022
rect 12893 23019 12959 23022
rect 19885 23082 19951 23085
rect 19885 23080 20178 23082
rect 19885 23024 19890 23080
rect 19946 23024 20178 23080
rect 19885 23022 20178 23024
rect 19885 23019 19951 23022
rect 3646 22880 4042 22881
rect 3646 22816 3652 22880
rect 3716 22816 3732 22880
rect 3796 22816 3812 22880
rect 3876 22816 3892 22880
rect 3956 22816 3972 22880
rect 4036 22816 4042 22880
rect 3646 22815 4042 22816
rect 7646 22880 8042 22881
rect 7646 22816 7652 22880
rect 7716 22816 7732 22880
rect 7796 22816 7812 22880
rect 7876 22816 7892 22880
rect 7956 22816 7972 22880
rect 8036 22816 8042 22880
rect 7646 22815 8042 22816
rect 11646 22880 12042 22881
rect 11646 22816 11652 22880
rect 11716 22816 11732 22880
rect 11796 22816 11812 22880
rect 11876 22816 11892 22880
rect 11956 22816 11972 22880
rect 12036 22816 12042 22880
rect 11646 22815 12042 22816
rect 15646 22880 16042 22881
rect 15646 22816 15652 22880
rect 15716 22816 15732 22880
rect 15796 22816 15812 22880
rect 15876 22816 15892 22880
rect 15956 22816 15972 22880
rect 16036 22816 16042 22880
rect 15646 22815 16042 22816
rect 19646 22880 20042 22881
rect 19646 22816 19652 22880
rect 19716 22816 19732 22880
rect 19796 22816 19812 22880
rect 19876 22816 19892 22880
rect 19956 22816 19972 22880
rect 20036 22816 20042 22880
rect 19646 22815 20042 22816
rect 19885 22674 19951 22677
rect 20118 22674 20178 23022
rect 23646 22880 24042 22881
rect 23646 22816 23652 22880
rect 23716 22816 23732 22880
rect 23796 22816 23812 22880
rect 23876 22816 23892 22880
rect 23956 22816 23972 22880
rect 24036 22816 24042 22880
rect 23646 22815 24042 22816
rect 19885 22672 20178 22674
rect 19885 22616 19890 22672
rect 19946 22616 20178 22672
rect 19885 22614 20178 22616
rect 19885 22611 19951 22614
rect 16573 22538 16639 22541
rect 17350 22538 17356 22540
rect 16573 22536 17356 22538
rect 16573 22480 16578 22536
rect 16634 22480 17356 22536
rect 16573 22478 17356 22480
rect 16573 22475 16639 22478
rect 17350 22476 17356 22478
rect 17420 22476 17426 22540
rect 26509 22538 26575 22541
rect 27171 22538 27971 22568
rect 26509 22536 27971 22538
rect 26509 22480 26514 22536
rect 26570 22480 27971 22536
rect 26509 22478 27971 22480
rect 26509 22475 26575 22478
rect 27171 22448 27971 22478
rect 2906 22336 3302 22337
rect 2906 22272 2912 22336
rect 2976 22272 2992 22336
rect 3056 22272 3072 22336
rect 3136 22272 3152 22336
rect 3216 22272 3232 22336
rect 3296 22272 3302 22336
rect 2906 22271 3302 22272
rect 6906 22336 7302 22337
rect 6906 22272 6912 22336
rect 6976 22272 6992 22336
rect 7056 22272 7072 22336
rect 7136 22272 7152 22336
rect 7216 22272 7232 22336
rect 7296 22272 7302 22336
rect 6906 22271 7302 22272
rect 10906 22336 11302 22337
rect 10906 22272 10912 22336
rect 10976 22272 10992 22336
rect 11056 22272 11072 22336
rect 11136 22272 11152 22336
rect 11216 22272 11232 22336
rect 11296 22272 11302 22336
rect 10906 22271 11302 22272
rect 14906 22336 15302 22337
rect 14906 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15072 22336
rect 15136 22272 15152 22336
rect 15216 22272 15232 22336
rect 15296 22272 15302 22336
rect 14906 22271 15302 22272
rect 18906 22336 19302 22337
rect 18906 22272 18912 22336
rect 18976 22272 18992 22336
rect 19056 22272 19072 22336
rect 19136 22272 19152 22336
rect 19216 22272 19232 22336
rect 19296 22272 19302 22336
rect 18906 22271 19302 22272
rect 22906 22336 23302 22337
rect 22906 22272 22912 22336
rect 22976 22272 22992 22336
rect 23056 22272 23072 22336
rect 23136 22272 23152 22336
rect 23216 22272 23232 22336
rect 23296 22272 23302 22336
rect 22906 22271 23302 22272
rect 5349 22132 5415 22133
rect 5349 22128 5396 22132
rect 5460 22130 5466 22132
rect 19885 22130 19951 22133
rect 20713 22130 20779 22133
rect 5349 22072 5354 22128
rect 5349 22068 5396 22072
rect 5460 22070 5506 22130
rect 19885 22128 20779 22130
rect 19885 22072 19890 22128
rect 19946 22072 20718 22128
rect 20774 22072 20779 22128
rect 19885 22070 20779 22072
rect 5460 22068 5466 22070
rect 5349 22067 5415 22068
rect 19885 22067 19951 22070
rect 20713 22067 20779 22070
rect 20529 21994 20595 21997
rect 24342 21994 24348 21996
rect 20529 21992 24348 21994
rect 20529 21936 20534 21992
rect 20590 21936 24348 21992
rect 20529 21934 24348 21936
rect 20529 21931 20595 21934
rect 24342 21932 24348 21934
rect 24412 21932 24418 21996
rect 3646 21792 4042 21793
rect 3646 21728 3652 21792
rect 3716 21728 3732 21792
rect 3796 21728 3812 21792
rect 3876 21728 3892 21792
rect 3956 21728 3972 21792
rect 4036 21728 4042 21792
rect 3646 21727 4042 21728
rect 7646 21792 8042 21793
rect 7646 21728 7652 21792
rect 7716 21728 7732 21792
rect 7796 21728 7812 21792
rect 7876 21728 7892 21792
rect 7956 21728 7972 21792
rect 8036 21728 8042 21792
rect 7646 21727 8042 21728
rect 11646 21792 12042 21793
rect 11646 21728 11652 21792
rect 11716 21728 11732 21792
rect 11796 21728 11812 21792
rect 11876 21728 11892 21792
rect 11956 21728 11972 21792
rect 12036 21728 12042 21792
rect 11646 21727 12042 21728
rect 15646 21792 16042 21793
rect 15646 21728 15652 21792
rect 15716 21728 15732 21792
rect 15796 21728 15812 21792
rect 15876 21728 15892 21792
rect 15956 21728 15972 21792
rect 16036 21728 16042 21792
rect 15646 21727 16042 21728
rect 19646 21792 20042 21793
rect 19646 21728 19652 21792
rect 19716 21728 19732 21792
rect 19796 21728 19812 21792
rect 19876 21728 19892 21792
rect 19956 21728 19972 21792
rect 20036 21728 20042 21792
rect 19646 21727 20042 21728
rect 23646 21792 24042 21793
rect 23646 21728 23652 21792
rect 23716 21728 23732 21792
rect 23796 21728 23812 21792
rect 23876 21728 23892 21792
rect 23956 21728 23972 21792
rect 24036 21728 24042 21792
rect 23646 21727 24042 21728
rect 2906 21248 3302 21249
rect 2906 21184 2912 21248
rect 2976 21184 2992 21248
rect 3056 21184 3072 21248
rect 3136 21184 3152 21248
rect 3216 21184 3232 21248
rect 3296 21184 3302 21248
rect 2906 21183 3302 21184
rect 6906 21248 7302 21249
rect 6906 21184 6912 21248
rect 6976 21184 6992 21248
rect 7056 21184 7072 21248
rect 7136 21184 7152 21248
rect 7216 21184 7232 21248
rect 7296 21184 7302 21248
rect 6906 21183 7302 21184
rect 10906 21248 11302 21249
rect 10906 21184 10912 21248
rect 10976 21184 10992 21248
rect 11056 21184 11072 21248
rect 11136 21184 11152 21248
rect 11216 21184 11232 21248
rect 11296 21184 11302 21248
rect 10906 21183 11302 21184
rect 14906 21248 15302 21249
rect 14906 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15072 21248
rect 15136 21184 15152 21248
rect 15216 21184 15232 21248
rect 15296 21184 15302 21248
rect 14906 21183 15302 21184
rect 18906 21248 19302 21249
rect 18906 21184 18912 21248
rect 18976 21184 18992 21248
rect 19056 21184 19072 21248
rect 19136 21184 19152 21248
rect 19216 21184 19232 21248
rect 19296 21184 19302 21248
rect 18906 21183 19302 21184
rect 22906 21248 23302 21249
rect 22906 21184 22912 21248
rect 22976 21184 22992 21248
rect 23056 21184 23072 21248
rect 23136 21184 23152 21248
rect 23216 21184 23232 21248
rect 23296 21184 23302 21248
rect 22906 21183 23302 21184
rect 19374 20844 19380 20908
rect 19444 20906 19450 20908
rect 19609 20906 19675 20909
rect 19444 20904 19675 20906
rect 19444 20848 19614 20904
rect 19670 20848 19675 20904
rect 19444 20846 19675 20848
rect 19444 20844 19450 20846
rect 19609 20843 19675 20846
rect 3646 20704 4042 20705
rect 3646 20640 3652 20704
rect 3716 20640 3732 20704
rect 3796 20640 3812 20704
rect 3876 20640 3892 20704
rect 3956 20640 3972 20704
rect 4036 20640 4042 20704
rect 3646 20639 4042 20640
rect 7646 20704 8042 20705
rect 7646 20640 7652 20704
rect 7716 20640 7732 20704
rect 7796 20640 7812 20704
rect 7876 20640 7892 20704
rect 7956 20640 7972 20704
rect 8036 20640 8042 20704
rect 7646 20639 8042 20640
rect 11646 20704 12042 20705
rect 11646 20640 11652 20704
rect 11716 20640 11732 20704
rect 11796 20640 11812 20704
rect 11876 20640 11892 20704
rect 11956 20640 11972 20704
rect 12036 20640 12042 20704
rect 11646 20639 12042 20640
rect 15646 20704 16042 20705
rect 15646 20640 15652 20704
rect 15716 20640 15732 20704
rect 15796 20640 15812 20704
rect 15876 20640 15892 20704
rect 15956 20640 15972 20704
rect 16036 20640 16042 20704
rect 15646 20639 16042 20640
rect 19646 20704 20042 20705
rect 19646 20640 19652 20704
rect 19716 20640 19732 20704
rect 19796 20640 19812 20704
rect 19876 20640 19892 20704
rect 19956 20640 19972 20704
rect 20036 20640 20042 20704
rect 19646 20639 20042 20640
rect 23646 20704 24042 20705
rect 23646 20640 23652 20704
rect 23716 20640 23732 20704
rect 23796 20640 23812 20704
rect 23876 20640 23892 20704
rect 23956 20640 23972 20704
rect 24036 20640 24042 20704
rect 23646 20639 24042 20640
rect 15469 20362 15535 20365
rect 18321 20364 18387 20365
rect 18270 20362 18276 20364
rect 15469 20360 18276 20362
rect 18340 20362 18387 20364
rect 18340 20360 18432 20362
rect 15469 20304 15474 20360
rect 15530 20304 18276 20360
rect 18382 20304 18432 20360
rect 15469 20302 18276 20304
rect 15469 20299 15535 20302
rect 18270 20300 18276 20302
rect 18340 20302 18432 20304
rect 18340 20300 18387 20302
rect 18321 20299 18387 20300
rect 2906 20160 3302 20161
rect 2906 20096 2912 20160
rect 2976 20096 2992 20160
rect 3056 20096 3072 20160
rect 3136 20096 3152 20160
rect 3216 20096 3232 20160
rect 3296 20096 3302 20160
rect 2906 20095 3302 20096
rect 6906 20160 7302 20161
rect 6906 20096 6912 20160
rect 6976 20096 6992 20160
rect 7056 20096 7072 20160
rect 7136 20096 7152 20160
rect 7216 20096 7232 20160
rect 7296 20096 7302 20160
rect 6906 20095 7302 20096
rect 10906 20160 11302 20161
rect 10906 20096 10912 20160
rect 10976 20096 10992 20160
rect 11056 20096 11072 20160
rect 11136 20096 11152 20160
rect 11216 20096 11232 20160
rect 11296 20096 11302 20160
rect 10906 20095 11302 20096
rect 14906 20160 15302 20161
rect 14906 20096 14912 20160
rect 14976 20096 14992 20160
rect 15056 20096 15072 20160
rect 15136 20096 15152 20160
rect 15216 20096 15232 20160
rect 15296 20096 15302 20160
rect 14906 20095 15302 20096
rect 18906 20160 19302 20161
rect 18906 20096 18912 20160
rect 18976 20096 18992 20160
rect 19056 20096 19072 20160
rect 19136 20096 19152 20160
rect 19216 20096 19232 20160
rect 19296 20096 19302 20160
rect 18906 20095 19302 20096
rect 22906 20160 23302 20161
rect 22906 20096 22912 20160
rect 22976 20096 22992 20160
rect 23056 20096 23072 20160
rect 23136 20096 23152 20160
rect 23216 20096 23232 20160
rect 23296 20096 23302 20160
rect 22906 20095 23302 20096
rect 3646 19616 4042 19617
rect 3646 19552 3652 19616
rect 3716 19552 3732 19616
rect 3796 19552 3812 19616
rect 3876 19552 3892 19616
rect 3956 19552 3972 19616
rect 4036 19552 4042 19616
rect 3646 19551 4042 19552
rect 7646 19616 8042 19617
rect 7646 19552 7652 19616
rect 7716 19552 7732 19616
rect 7796 19552 7812 19616
rect 7876 19552 7892 19616
rect 7956 19552 7972 19616
rect 8036 19552 8042 19616
rect 7646 19551 8042 19552
rect 11646 19616 12042 19617
rect 11646 19552 11652 19616
rect 11716 19552 11732 19616
rect 11796 19552 11812 19616
rect 11876 19552 11892 19616
rect 11956 19552 11972 19616
rect 12036 19552 12042 19616
rect 11646 19551 12042 19552
rect 15646 19616 16042 19617
rect 15646 19552 15652 19616
rect 15716 19552 15732 19616
rect 15796 19552 15812 19616
rect 15876 19552 15892 19616
rect 15956 19552 15972 19616
rect 16036 19552 16042 19616
rect 15646 19551 16042 19552
rect 19646 19616 20042 19617
rect 19646 19552 19652 19616
rect 19716 19552 19732 19616
rect 19796 19552 19812 19616
rect 19876 19552 19892 19616
rect 19956 19552 19972 19616
rect 20036 19552 20042 19616
rect 19646 19551 20042 19552
rect 23646 19616 24042 19617
rect 23646 19552 23652 19616
rect 23716 19552 23732 19616
rect 23796 19552 23812 19616
rect 23876 19552 23892 19616
rect 23956 19552 23972 19616
rect 24036 19552 24042 19616
rect 23646 19551 24042 19552
rect 5257 19412 5323 19413
rect 5206 19410 5212 19412
rect 5166 19350 5212 19410
rect 5276 19408 5323 19412
rect 5318 19352 5323 19408
rect 5206 19348 5212 19350
rect 5276 19348 5323 19352
rect 5257 19347 5323 19348
rect 5441 19410 5507 19413
rect 10409 19410 10475 19413
rect 5441 19408 10475 19410
rect 5441 19352 5446 19408
rect 5502 19352 10414 19408
rect 10470 19352 10475 19408
rect 5441 19350 10475 19352
rect 5441 19347 5507 19350
rect 10409 19347 10475 19350
rect 9990 19212 9996 19276
rect 10060 19274 10066 19276
rect 10225 19274 10291 19277
rect 10060 19272 10291 19274
rect 10060 19216 10230 19272
rect 10286 19216 10291 19272
rect 10060 19214 10291 19216
rect 10060 19212 10066 19214
rect 10225 19211 10291 19214
rect 2906 19072 3302 19073
rect 2906 19008 2912 19072
rect 2976 19008 2992 19072
rect 3056 19008 3072 19072
rect 3136 19008 3152 19072
rect 3216 19008 3232 19072
rect 3296 19008 3302 19072
rect 2906 19007 3302 19008
rect 6906 19072 7302 19073
rect 6906 19008 6912 19072
rect 6976 19008 6992 19072
rect 7056 19008 7072 19072
rect 7136 19008 7152 19072
rect 7216 19008 7232 19072
rect 7296 19008 7302 19072
rect 6906 19007 7302 19008
rect 10906 19072 11302 19073
rect 10906 19008 10912 19072
rect 10976 19008 10992 19072
rect 11056 19008 11072 19072
rect 11136 19008 11152 19072
rect 11216 19008 11232 19072
rect 11296 19008 11302 19072
rect 10906 19007 11302 19008
rect 14906 19072 15302 19073
rect 14906 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15072 19072
rect 15136 19008 15152 19072
rect 15216 19008 15232 19072
rect 15296 19008 15302 19072
rect 14906 19007 15302 19008
rect 18906 19072 19302 19073
rect 18906 19008 18912 19072
rect 18976 19008 18992 19072
rect 19056 19008 19072 19072
rect 19136 19008 19152 19072
rect 19216 19008 19232 19072
rect 19296 19008 19302 19072
rect 18906 19007 19302 19008
rect 22906 19072 23302 19073
rect 22906 19008 22912 19072
rect 22976 19008 22992 19072
rect 23056 19008 23072 19072
rect 23136 19008 23152 19072
rect 23216 19008 23232 19072
rect 23296 19008 23302 19072
rect 22906 19007 23302 19008
rect 9673 18866 9739 18869
rect 10317 18866 10383 18869
rect 9673 18864 10383 18866
rect 9673 18808 9678 18864
rect 9734 18808 10322 18864
rect 10378 18808 10383 18864
rect 9673 18806 10383 18808
rect 9673 18803 9739 18806
rect 10317 18803 10383 18806
rect 3646 18528 4042 18529
rect 3646 18464 3652 18528
rect 3716 18464 3732 18528
rect 3796 18464 3812 18528
rect 3876 18464 3892 18528
rect 3956 18464 3972 18528
rect 4036 18464 4042 18528
rect 3646 18463 4042 18464
rect 7646 18528 8042 18529
rect 7646 18464 7652 18528
rect 7716 18464 7732 18528
rect 7796 18464 7812 18528
rect 7876 18464 7892 18528
rect 7956 18464 7972 18528
rect 8036 18464 8042 18528
rect 7646 18463 8042 18464
rect 11646 18528 12042 18529
rect 11646 18464 11652 18528
rect 11716 18464 11732 18528
rect 11796 18464 11812 18528
rect 11876 18464 11892 18528
rect 11956 18464 11972 18528
rect 12036 18464 12042 18528
rect 11646 18463 12042 18464
rect 15646 18528 16042 18529
rect 15646 18464 15652 18528
rect 15716 18464 15732 18528
rect 15796 18464 15812 18528
rect 15876 18464 15892 18528
rect 15956 18464 15972 18528
rect 16036 18464 16042 18528
rect 15646 18463 16042 18464
rect 19646 18528 20042 18529
rect 19646 18464 19652 18528
rect 19716 18464 19732 18528
rect 19796 18464 19812 18528
rect 19876 18464 19892 18528
rect 19956 18464 19972 18528
rect 20036 18464 20042 18528
rect 19646 18463 20042 18464
rect 23646 18528 24042 18529
rect 23646 18464 23652 18528
rect 23716 18464 23732 18528
rect 23796 18464 23812 18528
rect 23876 18464 23892 18528
rect 23956 18464 23972 18528
rect 24036 18464 24042 18528
rect 23646 18463 24042 18464
rect 10409 18186 10475 18189
rect 14590 18186 14596 18188
rect 10409 18184 14596 18186
rect 10409 18128 10414 18184
rect 10470 18128 14596 18184
rect 10409 18126 14596 18128
rect 10409 18123 10475 18126
rect 14590 18124 14596 18126
rect 14660 18186 14666 18188
rect 17585 18186 17651 18189
rect 14660 18184 17651 18186
rect 14660 18128 17590 18184
rect 17646 18128 17651 18184
rect 14660 18126 17651 18128
rect 14660 18124 14666 18126
rect 17585 18123 17651 18126
rect 2906 17984 3302 17985
rect 2906 17920 2912 17984
rect 2976 17920 2992 17984
rect 3056 17920 3072 17984
rect 3136 17920 3152 17984
rect 3216 17920 3232 17984
rect 3296 17920 3302 17984
rect 2906 17919 3302 17920
rect 6906 17984 7302 17985
rect 6906 17920 6912 17984
rect 6976 17920 6992 17984
rect 7056 17920 7072 17984
rect 7136 17920 7152 17984
rect 7216 17920 7232 17984
rect 7296 17920 7302 17984
rect 6906 17919 7302 17920
rect 10906 17984 11302 17985
rect 10906 17920 10912 17984
rect 10976 17920 10992 17984
rect 11056 17920 11072 17984
rect 11136 17920 11152 17984
rect 11216 17920 11232 17984
rect 11296 17920 11302 17984
rect 10906 17919 11302 17920
rect 14906 17984 15302 17985
rect 14906 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15072 17984
rect 15136 17920 15152 17984
rect 15216 17920 15232 17984
rect 15296 17920 15302 17984
rect 14906 17919 15302 17920
rect 18906 17984 19302 17985
rect 18906 17920 18912 17984
rect 18976 17920 18992 17984
rect 19056 17920 19072 17984
rect 19136 17920 19152 17984
rect 19216 17920 19232 17984
rect 19296 17920 19302 17984
rect 18906 17919 19302 17920
rect 22906 17984 23302 17985
rect 22906 17920 22912 17984
rect 22976 17920 22992 17984
rect 23056 17920 23072 17984
rect 23136 17920 23152 17984
rect 23216 17920 23232 17984
rect 23296 17920 23302 17984
rect 22906 17919 23302 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 3646 17440 4042 17441
rect 3646 17376 3652 17440
rect 3716 17376 3732 17440
rect 3796 17376 3812 17440
rect 3876 17376 3892 17440
rect 3956 17376 3972 17440
rect 4036 17376 4042 17440
rect 3646 17375 4042 17376
rect 7646 17440 8042 17441
rect 7646 17376 7652 17440
rect 7716 17376 7732 17440
rect 7796 17376 7812 17440
rect 7876 17376 7892 17440
rect 7956 17376 7972 17440
rect 8036 17376 8042 17440
rect 7646 17375 8042 17376
rect 11646 17440 12042 17441
rect 11646 17376 11652 17440
rect 11716 17376 11732 17440
rect 11796 17376 11812 17440
rect 11876 17376 11892 17440
rect 11956 17376 11972 17440
rect 12036 17376 12042 17440
rect 11646 17375 12042 17376
rect 15646 17440 16042 17441
rect 15646 17376 15652 17440
rect 15716 17376 15732 17440
rect 15796 17376 15812 17440
rect 15876 17376 15892 17440
rect 15956 17376 15972 17440
rect 16036 17376 16042 17440
rect 15646 17375 16042 17376
rect 19646 17440 20042 17441
rect 19646 17376 19652 17440
rect 19716 17376 19732 17440
rect 19796 17376 19812 17440
rect 19876 17376 19892 17440
rect 19956 17376 19972 17440
rect 20036 17376 20042 17440
rect 19646 17375 20042 17376
rect 23646 17440 24042 17441
rect 23646 17376 23652 17440
rect 23716 17376 23732 17440
rect 23796 17376 23812 17440
rect 23876 17376 23892 17440
rect 23956 17376 23972 17440
rect 24036 17376 24042 17440
rect 23646 17375 24042 17376
rect 12893 17098 12959 17101
rect 18597 17098 18663 17101
rect 12893 17096 18663 17098
rect 12893 17040 12898 17096
rect 12954 17040 18602 17096
rect 18658 17040 18663 17096
rect 12893 17038 18663 17040
rect 12893 17035 12959 17038
rect 18597 17035 18663 17038
rect 2906 16896 3302 16897
rect 2906 16832 2912 16896
rect 2976 16832 2992 16896
rect 3056 16832 3072 16896
rect 3136 16832 3152 16896
rect 3216 16832 3232 16896
rect 3296 16832 3302 16896
rect 2906 16831 3302 16832
rect 6906 16896 7302 16897
rect 6906 16832 6912 16896
rect 6976 16832 6992 16896
rect 7056 16832 7072 16896
rect 7136 16832 7152 16896
rect 7216 16832 7232 16896
rect 7296 16832 7302 16896
rect 6906 16831 7302 16832
rect 10906 16896 11302 16897
rect 10906 16832 10912 16896
rect 10976 16832 10992 16896
rect 11056 16832 11072 16896
rect 11136 16832 11152 16896
rect 11216 16832 11232 16896
rect 11296 16832 11302 16896
rect 10906 16831 11302 16832
rect 14906 16896 15302 16897
rect 14906 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15072 16896
rect 15136 16832 15152 16896
rect 15216 16832 15232 16896
rect 15296 16832 15302 16896
rect 14906 16831 15302 16832
rect 18906 16896 19302 16897
rect 18906 16832 18912 16896
rect 18976 16832 18992 16896
rect 19056 16832 19072 16896
rect 19136 16832 19152 16896
rect 19216 16832 19232 16896
rect 19296 16832 19302 16896
rect 18906 16831 19302 16832
rect 22906 16896 23302 16897
rect 22906 16832 22912 16896
rect 22976 16832 22992 16896
rect 23056 16832 23072 16896
rect 23136 16832 23152 16896
rect 23216 16832 23232 16896
rect 23296 16832 23302 16896
rect 22906 16831 23302 16832
rect 15561 16692 15627 16693
rect 15510 16690 15516 16692
rect 15470 16630 15516 16690
rect 15580 16688 15627 16692
rect 15622 16632 15627 16688
rect 15510 16628 15516 16630
rect 15580 16628 15627 16632
rect 15561 16627 15627 16628
rect 13629 16554 13695 16557
rect 18965 16554 19031 16557
rect 13629 16552 19031 16554
rect 13629 16496 13634 16552
rect 13690 16496 18970 16552
rect 19026 16496 19031 16552
rect 13629 16494 19031 16496
rect 13629 16491 13695 16494
rect 18965 16491 19031 16494
rect 3646 16352 4042 16353
rect 3646 16288 3652 16352
rect 3716 16288 3732 16352
rect 3796 16288 3812 16352
rect 3876 16288 3892 16352
rect 3956 16288 3972 16352
rect 4036 16288 4042 16352
rect 3646 16287 4042 16288
rect 7646 16352 8042 16353
rect 7646 16288 7652 16352
rect 7716 16288 7732 16352
rect 7796 16288 7812 16352
rect 7876 16288 7892 16352
rect 7956 16288 7972 16352
rect 8036 16288 8042 16352
rect 7646 16287 8042 16288
rect 11646 16352 12042 16353
rect 11646 16288 11652 16352
rect 11716 16288 11732 16352
rect 11796 16288 11812 16352
rect 11876 16288 11892 16352
rect 11956 16288 11972 16352
rect 12036 16288 12042 16352
rect 11646 16287 12042 16288
rect 15646 16352 16042 16353
rect 15646 16288 15652 16352
rect 15716 16288 15732 16352
rect 15796 16288 15812 16352
rect 15876 16288 15892 16352
rect 15956 16288 15972 16352
rect 16036 16288 16042 16352
rect 15646 16287 16042 16288
rect 19646 16352 20042 16353
rect 19646 16288 19652 16352
rect 19716 16288 19732 16352
rect 19796 16288 19812 16352
rect 19876 16288 19892 16352
rect 19956 16288 19972 16352
rect 20036 16288 20042 16352
rect 19646 16287 20042 16288
rect 23646 16352 24042 16353
rect 23646 16288 23652 16352
rect 23716 16288 23732 16352
rect 23796 16288 23812 16352
rect 23876 16288 23892 16352
rect 23956 16288 23972 16352
rect 24036 16288 24042 16352
rect 23646 16287 24042 16288
rect 17769 16282 17835 16285
rect 18638 16282 18644 16284
rect 17769 16280 18644 16282
rect 17769 16224 17774 16280
rect 17830 16224 18644 16280
rect 17769 16222 18644 16224
rect 17769 16219 17835 16222
rect 18638 16220 18644 16222
rect 18708 16282 18714 16284
rect 18781 16282 18847 16285
rect 19333 16284 19399 16285
rect 19333 16282 19380 16284
rect 18708 16280 18847 16282
rect 18708 16224 18786 16280
rect 18842 16224 18847 16280
rect 18708 16222 18847 16224
rect 19288 16280 19380 16282
rect 19288 16224 19338 16280
rect 19288 16222 19380 16224
rect 18708 16220 18714 16222
rect 18781 16219 18847 16222
rect 19333 16220 19380 16222
rect 19444 16220 19450 16284
rect 19333 16219 19399 16220
rect 14590 16084 14596 16148
rect 14660 16146 14666 16148
rect 21817 16146 21883 16149
rect 14660 16144 21883 16146
rect 14660 16088 21822 16144
rect 21878 16088 21883 16144
rect 14660 16086 21883 16088
rect 14660 16084 14666 16086
rect 21817 16083 21883 16086
rect 10869 16010 10935 16013
rect 16573 16010 16639 16013
rect 10869 16008 16639 16010
rect 10869 15952 10874 16008
rect 10930 15952 16578 16008
rect 16634 15952 16639 16008
rect 10869 15950 16639 15952
rect 10869 15947 10935 15950
rect 16573 15947 16639 15950
rect 2906 15808 3302 15809
rect 2906 15744 2912 15808
rect 2976 15744 2992 15808
rect 3056 15744 3072 15808
rect 3136 15744 3152 15808
rect 3216 15744 3232 15808
rect 3296 15744 3302 15808
rect 2906 15743 3302 15744
rect 6906 15808 7302 15809
rect 6906 15744 6912 15808
rect 6976 15744 6992 15808
rect 7056 15744 7072 15808
rect 7136 15744 7152 15808
rect 7216 15744 7232 15808
rect 7296 15744 7302 15808
rect 6906 15743 7302 15744
rect 10906 15808 11302 15809
rect 10906 15744 10912 15808
rect 10976 15744 10992 15808
rect 11056 15744 11072 15808
rect 11136 15744 11152 15808
rect 11216 15744 11232 15808
rect 11296 15744 11302 15808
rect 10906 15743 11302 15744
rect 14906 15808 15302 15809
rect 14906 15744 14912 15808
rect 14976 15744 14992 15808
rect 15056 15744 15072 15808
rect 15136 15744 15152 15808
rect 15216 15744 15232 15808
rect 15296 15744 15302 15808
rect 14906 15743 15302 15744
rect 18906 15808 19302 15809
rect 18906 15744 18912 15808
rect 18976 15744 18992 15808
rect 19056 15744 19072 15808
rect 19136 15744 19152 15808
rect 19216 15744 19232 15808
rect 19296 15744 19302 15808
rect 18906 15743 19302 15744
rect 22906 15808 23302 15809
rect 22906 15744 22912 15808
rect 22976 15744 22992 15808
rect 23056 15744 23072 15808
rect 23136 15744 23152 15808
rect 23216 15744 23232 15808
rect 23296 15744 23302 15808
rect 22906 15743 23302 15744
rect 10501 15466 10567 15469
rect 18229 15466 18295 15469
rect 10501 15464 18295 15466
rect 10501 15408 10506 15464
rect 10562 15408 18234 15464
rect 18290 15408 18295 15464
rect 10501 15406 18295 15408
rect 10501 15403 10567 15406
rect 18229 15403 18295 15406
rect 3646 15264 4042 15265
rect 3646 15200 3652 15264
rect 3716 15200 3732 15264
rect 3796 15200 3812 15264
rect 3876 15200 3892 15264
rect 3956 15200 3972 15264
rect 4036 15200 4042 15264
rect 3646 15199 4042 15200
rect 7646 15264 8042 15265
rect 7646 15200 7652 15264
rect 7716 15200 7732 15264
rect 7796 15200 7812 15264
rect 7876 15200 7892 15264
rect 7956 15200 7972 15264
rect 8036 15200 8042 15264
rect 7646 15199 8042 15200
rect 11646 15264 12042 15265
rect 11646 15200 11652 15264
rect 11716 15200 11732 15264
rect 11796 15200 11812 15264
rect 11876 15200 11892 15264
rect 11956 15200 11972 15264
rect 12036 15200 12042 15264
rect 11646 15199 12042 15200
rect 15646 15264 16042 15265
rect 15646 15200 15652 15264
rect 15716 15200 15732 15264
rect 15796 15200 15812 15264
rect 15876 15200 15892 15264
rect 15956 15200 15972 15264
rect 16036 15200 16042 15264
rect 15646 15199 16042 15200
rect 19646 15264 20042 15265
rect 19646 15200 19652 15264
rect 19716 15200 19732 15264
rect 19796 15200 19812 15264
rect 19876 15200 19892 15264
rect 19956 15200 19972 15264
rect 20036 15200 20042 15264
rect 19646 15199 20042 15200
rect 23646 15264 24042 15265
rect 23646 15200 23652 15264
rect 23716 15200 23732 15264
rect 23796 15200 23812 15264
rect 23876 15200 23892 15264
rect 23956 15200 23972 15264
rect 24036 15200 24042 15264
rect 23646 15199 24042 15200
rect 9121 15194 9187 15197
rect 11053 15194 11119 15197
rect 9121 15192 11119 15194
rect 9121 15136 9126 15192
rect 9182 15136 11058 15192
rect 11114 15136 11119 15192
rect 9121 15134 11119 15136
rect 9121 15131 9187 15134
rect 11053 15131 11119 15134
rect 3417 15058 3483 15061
rect 13997 15058 14063 15061
rect 3417 15056 14063 15058
rect 3417 15000 3422 15056
rect 3478 15000 14002 15056
rect 14058 15000 14063 15056
rect 3417 14998 14063 15000
rect 3417 14995 3483 14998
rect 13997 14995 14063 14998
rect 7741 14922 7807 14925
rect 9029 14922 9095 14925
rect 7741 14920 9095 14922
rect 7741 14864 7746 14920
rect 7802 14864 9034 14920
rect 9090 14864 9095 14920
rect 7741 14862 9095 14864
rect 7741 14859 7807 14862
rect 9029 14859 9095 14862
rect 2906 14720 3302 14721
rect 2906 14656 2912 14720
rect 2976 14656 2992 14720
rect 3056 14656 3072 14720
rect 3136 14656 3152 14720
rect 3216 14656 3232 14720
rect 3296 14656 3302 14720
rect 2906 14655 3302 14656
rect 6906 14720 7302 14721
rect 6906 14656 6912 14720
rect 6976 14656 6992 14720
rect 7056 14656 7072 14720
rect 7136 14656 7152 14720
rect 7216 14656 7232 14720
rect 7296 14656 7302 14720
rect 6906 14655 7302 14656
rect 10906 14720 11302 14721
rect 10906 14656 10912 14720
rect 10976 14656 10992 14720
rect 11056 14656 11072 14720
rect 11136 14656 11152 14720
rect 11216 14656 11232 14720
rect 11296 14656 11302 14720
rect 10906 14655 11302 14656
rect 14906 14720 15302 14721
rect 14906 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15072 14720
rect 15136 14656 15152 14720
rect 15216 14656 15232 14720
rect 15296 14656 15302 14720
rect 14906 14655 15302 14656
rect 18906 14720 19302 14721
rect 18906 14656 18912 14720
rect 18976 14656 18992 14720
rect 19056 14656 19072 14720
rect 19136 14656 19152 14720
rect 19216 14656 19232 14720
rect 19296 14656 19302 14720
rect 18906 14655 19302 14656
rect 22906 14720 23302 14721
rect 22906 14656 22912 14720
rect 22976 14656 22992 14720
rect 23056 14656 23072 14720
rect 23136 14656 23152 14720
rect 23216 14656 23232 14720
rect 23296 14656 23302 14720
rect 22906 14655 23302 14656
rect 14590 14452 14596 14516
rect 14660 14514 14666 14516
rect 14825 14514 14891 14517
rect 14660 14512 14891 14514
rect 14660 14456 14830 14512
rect 14886 14456 14891 14512
rect 14660 14454 14891 14456
rect 14660 14452 14666 14454
rect 14825 14451 14891 14454
rect 15510 14452 15516 14516
rect 15580 14514 15586 14516
rect 15745 14514 15811 14517
rect 15580 14512 15811 14514
rect 15580 14456 15750 14512
rect 15806 14456 15811 14512
rect 15580 14454 15811 14456
rect 15580 14452 15586 14454
rect 13445 14378 13511 14381
rect 15518 14378 15578 14452
rect 15745 14451 15811 14454
rect 13445 14376 15578 14378
rect 13445 14320 13450 14376
rect 13506 14320 15578 14376
rect 13445 14318 15578 14320
rect 13445 14315 13511 14318
rect 18270 14316 18276 14380
rect 18340 14378 18346 14380
rect 18689 14378 18755 14381
rect 18340 14376 18755 14378
rect 18340 14320 18694 14376
rect 18750 14320 18755 14376
rect 18340 14318 18755 14320
rect 18340 14316 18346 14318
rect 18689 14315 18755 14318
rect 3646 14176 4042 14177
rect 3646 14112 3652 14176
rect 3716 14112 3732 14176
rect 3796 14112 3812 14176
rect 3876 14112 3892 14176
rect 3956 14112 3972 14176
rect 4036 14112 4042 14176
rect 3646 14111 4042 14112
rect 7646 14176 8042 14177
rect 7646 14112 7652 14176
rect 7716 14112 7732 14176
rect 7796 14112 7812 14176
rect 7876 14112 7892 14176
rect 7956 14112 7972 14176
rect 8036 14112 8042 14176
rect 7646 14111 8042 14112
rect 11646 14176 12042 14177
rect 11646 14112 11652 14176
rect 11716 14112 11732 14176
rect 11796 14112 11812 14176
rect 11876 14112 11892 14176
rect 11956 14112 11972 14176
rect 12036 14112 12042 14176
rect 11646 14111 12042 14112
rect 15646 14176 16042 14177
rect 15646 14112 15652 14176
rect 15716 14112 15732 14176
rect 15796 14112 15812 14176
rect 15876 14112 15892 14176
rect 15956 14112 15972 14176
rect 16036 14112 16042 14176
rect 15646 14111 16042 14112
rect 19646 14176 20042 14177
rect 19646 14112 19652 14176
rect 19716 14112 19732 14176
rect 19796 14112 19812 14176
rect 19876 14112 19892 14176
rect 19956 14112 19972 14176
rect 20036 14112 20042 14176
rect 19646 14111 20042 14112
rect 23646 14176 24042 14177
rect 23646 14112 23652 14176
rect 23716 14112 23732 14176
rect 23796 14112 23812 14176
rect 23876 14112 23892 14176
rect 23956 14112 23972 14176
rect 24036 14112 24042 14176
rect 23646 14111 24042 14112
rect 25957 13698 26023 13701
rect 27171 13698 27971 13728
rect 25957 13696 27971 13698
rect 25957 13640 25962 13696
rect 26018 13640 27971 13696
rect 25957 13638 27971 13640
rect 25957 13635 26023 13638
rect 2906 13632 3302 13633
rect 2906 13568 2912 13632
rect 2976 13568 2992 13632
rect 3056 13568 3072 13632
rect 3136 13568 3152 13632
rect 3216 13568 3232 13632
rect 3296 13568 3302 13632
rect 2906 13567 3302 13568
rect 6906 13632 7302 13633
rect 6906 13568 6912 13632
rect 6976 13568 6992 13632
rect 7056 13568 7072 13632
rect 7136 13568 7152 13632
rect 7216 13568 7232 13632
rect 7296 13568 7302 13632
rect 6906 13567 7302 13568
rect 10906 13632 11302 13633
rect 10906 13568 10912 13632
rect 10976 13568 10992 13632
rect 11056 13568 11072 13632
rect 11136 13568 11152 13632
rect 11216 13568 11232 13632
rect 11296 13568 11302 13632
rect 10906 13567 11302 13568
rect 14906 13632 15302 13633
rect 14906 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15072 13632
rect 15136 13568 15152 13632
rect 15216 13568 15232 13632
rect 15296 13568 15302 13632
rect 14906 13567 15302 13568
rect 18906 13632 19302 13633
rect 18906 13568 18912 13632
rect 18976 13568 18992 13632
rect 19056 13568 19072 13632
rect 19136 13568 19152 13632
rect 19216 13568 19232 13632
rect 19296 13568 19302 13632
rect 18906 13567 19302 13568
rect 22906 13632 23302 13633
rect 22906 13568 22912 13632
rect 22976 13568 22992 13632
rect 23056 13568 23072 13632
rect 23136 13568 23152 13632
rect 23216 13568 23232 13632
rect 23296 13568 23302 13632
rect 27171 13608 27971 13638
rect 22906 13567 23302 13568
rect 18413 13428 18479 13429
rect 18413 13424 18460 13428
rect 18524 13426 18530 13428
rect 18413 13368 18418 13424
rect 18413 13364 18460 13368
rect 18524 13366 18570 13426
rect 18524 13364 18530 13366
rect 18413 13363 18479 13364
rect 3646 13088 4042 13089
rect 0 13018 800 13048
rect 3646 13024 3652 13088
rect 3716 13024 3732 13088
rect 3796 13024 3812 13088
rect 3876 13024 3892 13088
rect 3956 13024 3972 13088
rect 4036 13024 4042 13088
rect 3646 13023 4042 13024
rect 7646 13088 8042 13089
rect 7646 13024 7652 13088
rect 7716 13024 7732 13088
rect 7796 13024 7812 13088
rect 7876 13024 7892 13088
rect 7956 13024 7972 13088
rect 8036 13024 8042 13088
rect 7646 13023 8042 13024
rect 11646 13088 12042 13089
rect 11646 13024 11652 13088
rect 11716 13024 11732 13088
rect 11796 13024 11812 13088
rect 11876 13024 11892 13088
rect 11956 13024 11972 13088
rect 12036 13024 12042 13088
rect 11646 13023 12042 13024
rect 15646 13088 16042 13089
rect 15646 13024 15652 13088
rect 15716 13024 15732 13088
rect 15796 13024 15812 13088
rect 15876 13024 15892 13088
rect 15956 13024 15972 13088
rect 16036 13024 16042 13088
rect 15646 13023 16042 13024
rect 19646 13088 20042 13089
rect 19646 13024 19652 13088
rect 19716 13024 19732 13088
rect 19796 13024 19812 13088
rect 19876 13024 19892 13088
rect 19956 13024 19972 13088
rect 20036 13024 20042 13088
rect 19646 13023 20042 13024
rect 23646 13088 24042 13089
rect 23646 13024 23652 13088
rect 23716 13024 23732 13088
rect 23796 13024 23812 13088
rect 23876 13024 23892 13088
rect 23956 13024 23972 13088
rect 24036 13024 24042 13088
rect 23646 13023 24042 13024
rect 0 12928 858 13018
rect 798 12885 858 12928
rect 798 12880 907 12885
rect 798 12824 846 12880
rect 902 12824 907 12880
rect 798 12822 907 12824
rect 841 12819 907 12822
rect 4705 12882 4771 12885
rect 5257 12884 5323 12885
rect 4705 12880 5090 12882
rect 4705 12824 4710 12880
rect 4766 12824 5090 12880
rect 4705 12822 5090 12824
rect 4705 12819 4771 12822
rect 5030 12746 5090 12822
rect 5206 12820 5212 12884
rect 5276 12882 5323 12884
rect 5276 12880 5368 12882
rect 5318 12824 5368 12880
rect 5276 12822 5368 12824
rect 5276 12820 5323 12822
rect 5257 12819 5323 12820
rect 5030 12686 5412 12746
rect 2906 12544 3302 12545
rect 2906 12480 2912 12544
rect 2976 12480 2992 12544
rect 3056 12480 3072 12544
rect 3136 12480 3152 12544
rect 3216 12480 3232 12544
rect 3296 12480 3302 12544
rect 2906 12479 3302 12480
rect 5352 12477 5412 12686
rect 6906 12544 7302 12545
rect 6906 12480 6912 12544
rect 6976 12480 6992 12544
rect 7056 12480 7072 12544
rect 7136 12480 7152 12544
rect 7216 12480 7232 12544
rect 7296 12480 7302 12544
rect 6906 12479 7302 12480
rect 10906 12544 11302 12545
rect 10906 12480 10912 12544
rect 10976 12480 10992 12544
rect 11056 12480 11072 12544
rect 11136 12480 11152 12544
rect 11216 12480 11232 12544
rect 11296 12480 11302 12544
rect 10906 12479 11302 12480
rect 14906 12544 15302 12545
rect 14906 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15072 12544
rect 15136 12480 15152 12544
rect 15216 12480 15232 12544
rect 15296 12480 15302 12544
rect 14906 12479 15302 12480
rect 18906 12544 19302 12545
rect 18906 12480 18912 12544
rect 18976 12480 18992 12544
rect 19056 12480 19072 12544
rect 19136 12480 19152 12544
rect 19216 12480 19232 12544
rect 19296 12480 19302 12544
rect 18906 12479 19302 12480
rect 22906 12544 23302 12545
rect 22906 12480 22912 12544
rect 22976 12480 22992 12544
rect 23056 12480 23072 12544
rect 23136 12480 23152 12544
rect 23216 12480 23232 12544
rect 23296 12480 23302 12544
rect 22906 12479 23302 12480
rect 5349 12472 5415 12477
rect 5349 12416 5354 12472
rect 5410 12416 5415 12472
rect 5349 12411 5415 12416
rect 3646 12000 4042 12001
rect 3646 11936 3652 12000
rect 3716 11936 3732 12000
rect 3796 11936 3812 12000
rect 3876 11936 3892 12000
rect 3956 11936 3972 12000
rect 4036 11936 4042 12000
rect 3646 11935 4042 11936
rect 7646 12000 8042 12001
rect 7646 11936 7652 12000
rect 7716 11936 7732 12000
rect 7796 11936 7812 12000
rect 7876 11936 7892 12000
rect 7956 11936 7972 12000
rect 8036 11936 8042 12000
rect 7646 11935 8042 11936
rect 11646 12000 12042 12001
rect 11646 11936 11652 12000
rect 11716 11936 11732 12000
rect 11796 11936 11812 12000
rect 11876 11936 11892 12000
rect 11956 11936 11972 12000
rect 12036 11936 12042 12000
rect 11646 11935 12042 11936
rect 15646 12000 16042 12001
rect 15646 11936 15652 12000
rect 15716 11936 15732 12000
rect 15796 11936 15812 12000
rect 15876 11936 15892 12000
rect 15956 11936 15972 12000
rect 16036 11936 16042 12000
rect 15646 11935 16042 11936
rect 19646 12000 20042 12001
rect 19646 11936 19652 12000
rect 19716 11936 19732 12000
rect 19796 11936 19812 12000
rect 19876 11936 19892 12000
rect 19956 11936 19972 12000
rect 20036 11936 20042 12000
rect 19646 11935 20042 11936
rect 23646 12000 24042 12001
rect 23646 11936 23652 12000
rect 23716 11936 23732 12000
rect 23796 11936 23812 12000
rect 23876 11936 23892 12000
rect 23956 11936 23972 12000
rect 24036 11936 24042 12000
rect 23646 11935 24042 11936
rect 5390 11732 5396 11796
rect 5460 11794 5466 11796
rect 9121 11794 9187 11797
rect 5460 11792 9187 11794
rect 5460 11736 9126 11792
rect 9182 11736 9187 11792
rect 5460 11734 9187 11736
rect 5460 11732 5466 11734
rect 9121 11731 9187 11734
rect 3693 11658 3759 11661
rect 9990 11658 9996 11660
rect 3693 11656 9996 11658
rect 3693 11600 3698 11656
rect 3754 11600 9996 11656
rect 3693 11598 9996 11600
rect 3693 11595 3759 11598
rect 9990 11596 9996 11598
rect 10060 11596 10066 11660
rect 2906 11456 3302 11457
rect 2906 11392 2912 11456
rect 2976 11392 2992 11456
rect 3056 11392 3072 11456
rect 3136 11392 3152 11456
rect 3216 11392 3232 11456
rect 3296 11392 3302 11456
rect 2906 11391 3302 11392
rect 6906 11456 7302 11457
rect 6906 11392 6912 11456
rect 6976 11392 6992 11456
rect 7056 11392 7072 11456
rect 7136 11392 7152 11456
rect 7216 11392 7232 11456
rect 7296 11392 7302 11456
rect 6906 11391 7302 11392
rect 10906 11456 11302 11457
rect 10906 11392 10912 11456
rect 10976 11392 10992 11456
rect 11056 11392 11072 11456
rect 11136 11392 11152 11456
rect 11216 11392 11232 11456
rect 11296 11392 11302 11456
rect 10906 11391 11302 11392
rect 14906 11456 15302 11457
rect 14906 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15072 11456
rect 15136 11392 15152 11456
rect 15216 11392 15232 11456
rect 15296 11392 15302 11456
rect 14906 11391 15302 11392
rect 18906 11456 19302 11457
rect 18906 11392 18912 11456
rect 18976 11392 18992 11456
rect 19056 11392 19072 11456
rect 19136 11392 19152 11456
rect 19216 11392 19232 11456
rect 19296 11392 19302 11456
rect 18906 11391 19302 11392
rect 22906 11456 23302 11457
rect 22906 11392 22912 11456
rect 22976 11392 22992 11456
rect 23056 11392 23072 11456
rect 23136 11392 23152 11456
rect 23216 11392 23232 11456
rect 23296 11392 23302 11456
rect 22906 11391 23302 11392
rect 3646 10912 4042 10913
rect 3646 10848 3652 10912
rect 3716 10848 3732 10912
rect 3796 10848 3812 10912
rect 3876 10848 3892 10912
rect 3956 10848 3972 10912
rect 4036 10848 4042 10912
rect 3646 10847 4042 10848
rect 7646 10912 8042 10913
rect 7646 10848 7652 10912
rect 7716 10848 7732 10912
rect 7796 10848 7812 10912
rect 7876 10848 7892 10912
rect 7956 10848 7972 10912
rect 8036 10848 8042 10912
rect 7646 10847 8042 10848
rect 11646 10912 12042 10913
rect 11646 10848 11652 10912
rect 11716 10848 11732 10912
rect 11796 10848 11812 10912
rect 11876 10848 11892 10912
rect 11956 10848 11972 10912
rect 12036 10848 12042 10912
rect 11646 10847 12042 10848
rect 15646 10912 16042 10913
rect 15646 10848 15652 10912
rect 15716 10848 15732 10912
rect 15796 10848 15812 10912
rect 15876 10848 15892 10912
rect 15956 10848 15972 10912
rect 16036 10848 16042 10912
rect 15646 10847 16042 10848
rect 19646 10912 20042 10913
rect 19646 10848 19652 10912
rect 19716 10848 19732 10912
rect 19796 10848 19812 10912
rect 19876 10848 19892 10912
rect 19956 10848 19972 10912
rect 20036 10848 20042 10912
rect 19646 10847 20042 10848
rect 23646 10912 24042 10913
rect 23646 10848 23652 10912
rect 23716 10848 23732 10912
rect 23796 10848 23812 10912
rect 23876 10848 23892 10912
rect 23956 10848 23972 10912
rect 24036 10848 24042 10912
rect 23646 10847 24042 10848
rect 10041 10842 10107 10845
rect 10174 10842 10180 10844
rect 10041 10840 10180 10842
rect 10041 10784 10046 10840
rect 10102 10784 10180 10840
rect 10041 10782 10180 10784
rect 10041 10779 10107 10782
rect 10174 10780 10180 10782
rect 10244 10780 10250 10844
rect 17309 10708 17375 10709
rect 17309 10706 17356 10708
rect 17264 10704 17356 10706
rect 17264 10648 17314 10704
rect 17264 10646 17356 10648
rect 17309 10644 17356 10646
rect 17420 10644 17426 10708
rect 17309 10643 17375 10644
rect 8109 10570 8175 10573
rect 8293 10570 8359 10573
rect 8109 10568 8359 10570
rect 8109 10512 8114 10568
rect 8170 10512 8298 10568
rect 8354 10512 8359 10568
rect 8109 10510 8359 10512
rect 8109 10507 8175 10510
rect 8293 10507 8359 10510
rect 2906 10368 3302 10369
rect 2906 10304 2912 10368
rect 2976 10304 2992 10368
rect 3056 10304 3072 10368
rect 3136 10304 3152 10368
rect 3216 10304 3232 10368
rect 3296 10304 3302 10368
rect 2906 10303 3302 10304
rect 6906 10368 7302 10369
rect 6906 10304 6912 10368
rect 6976 10304 6992 10368
rect 7056 10304 7072 10368
rect 7136 10304 7152 10368
rect 7216 10304 7232 10368
rect 7296 10304 7302 10368
rect 6906 10303 7302 10304
rect 10906 10368 11302 10369
rect 10906 10304 10912 10368
rect 10976 10304 10992 10368
rect 11056 10304 11072 10368
rect 11136 10304 11152 10368
rect 11216 10304 11232 10368
rect 11296 10304 11302 10368
rect 10906 10303 11302 10304
rect 14906 10368 15302 10369
rect 14906 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15072 10368
rect 15136 10304 15152 10368
rect 15216 10304 15232 10368
rect 15296 10304 15302 10368
rect 14906 10303 15302 10304
rect 18906 10368 19302 10369
rect 18906 10304 18912 10368
rect 18976 10304 18992 10368
rect 19056 10304 19072 10368
rect 19136 10304 19152 10368
rect 19216 10304 19232 10368
rect 19296 10304 19302 10368
rect 18906 10303 19302 10304
rect 22906 10368 23302 10369
rect 22906 10304 22912 10368
rect 22976 10304 22992 10368
rect 23056 10304 23072 10368
rect 23136 10304 23152 10368
rect 23216 10304 23232 10368
rect 23296 10304 23302 10368
rect 22906 10303 23302 10304
rect 7557 10298 7623 10301
rect 9489 10298 9555 10301
rect 17493 10300 17559 10301
rect 17493 10298 17540 10300
rect 7557 10296 9555 10298
rect 7557 10240 7562 10296
rect 7618 10240 9494 10296
rect 9550 10240 9555 10296
rect 7557 10238 9555 10240
rect 17448 10296 17540 10298
rect 17448 10240 17498 10296
rect 17448 10238 17540 10240
rect 7557 10235 7623 10238
rect 9489 10235 9555 10238
rect 17493 10236 17540 10238
rect 17604 10236 17610 10300
rect 18270 10236 18276 10300
rect 18340 10298 18346 10300
rect 18597 10298 18663 10301
rect 18340 10296 18663 10298
rect 18340 10240 18602 10296
rect 18658 10240 18663 10296
rect 18340 10238 18663 10240
rect 18340 10236 18346 10238
rect 17493 10235 17559 10236
rect 18597 10235 18663 10238
rect 7097 10162 7163 10165
rect 9029 10162 9095 10165
rect 7097 10160 9095 10162
rect 7097 10104 7102 10160
rect 7158 10104 9034 10160
rect 9090 10104 9095 10160
rect 7097 10102 9095 10104
rect 7097 10099 7163 10102
rect 9029 10099 9095 10102
rect 2681 10026 2747 10029
rect 3509 10026 3575 10029
rect 8477 10026 8543 10029
rect 9581 10026 9647 10029
rect 2681 10024 9647 10026
rect 2681 9968 2686 10024
rect 2742 9968 3514 10024
rect 3570 9968 8482 10024
rect 8538 9968 9586 10024
rect 9642 9968 9647 10024
rect 2681 9966 9647 9968
rect 2681 9963 2747 9966
rect 3509 9963 3575 9966
rect 8477 9963 8543 9966
rect 9581 9963 9647 9966
rect 14273 10026 14339 10029
rect 17585 10026 17651 10029
rect 14273 10024 17651 10026
rect 14273 9968 14278 10024
rect 14334 9968 17590 10024
rect 17646 9968 17651 10024
rect 14273 9966 17651 9968
rect 14273 9963 14339 9966
rect 17585 9963 17651 9966
rect 3646 9824 4042 9825
rect 3646 9760 3652 9824
rect 3716 9760 3732 9824
rect 3796 9760 3812 9824
rect 3876 9760 3892 9824
rect 3956 9760 3972 9824
rect 4036 9760 4042 9824
rect 3646 9759 4042 9760
rect 7646 9824 8042 9825
rect 7646 9760 7652 9824
rect 7716 9760 7732 9824
rect 7796 9760 7812 9824
rect 7876 9760 7892 9824
rect 7956 9760 7972 9824
rect 8036 9760 8042 9824
rect 7646 9759 8042 9760
rect 11646 9824 12042 9825
rect 11646 9760 11652 9824
rect 11716 9760 11732 9824
rect 11796 9760 11812 9824
rect 11876 9760 11892 9824
rect 11956 9760 11972 9824
rect 12036 9760 12042 9824
rect 11646 9759 12042 9760
rect 15646 9824 16042 9825
rect 15646 9760 15652 9824
rect 15716 9760 15732 9824
rect 15796 9760 15812 9824
rect 15876 9760 15892 9824
rect 15956 9760 15972 9824
rect 16036 9760 16042 9824
rect 15646 9759 16042 9760
rect 19646 9824 20042 9825
rect 19646 9760 19652 9824
rect 19716 9760 19732 9824
rect 19796 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20042 9824
rect 19646 9759 20042 9760
rect 23646 9824 24042 9825
rect 23646 9760 23652 9824
rect 23716 9760 23732 9824
rect 23796 9760 23812 9824
rect 23876 9760 23892 9824
rect 23956 9760 23972 9824
rect 24036 9760 24042 9824
rect 23646 9759 24042 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 26141 9618 26207 9621
rect 27171 9618 27971 9648
rect 26141 9616 27971 9618
rect 26141 9560 26146 9616
rect 26202 9560 27971 9616
rect 26141 9558 27971 9560
rect 26141 9555 26207 9558
rect 27171 9528 27971 9558
rect 2906 9280 3302 9281
rect 2906 9216 2912 9280
rect 2976 9216 2992 9280
rect 3056 9216 3072 9280
rect 3136 9216 3152 9280
rect 3216 9216 3232 9280
rect 3296 9216 3302 9280
rect 2906 9215 3302 9216
rect 6906 9280 7302 9281
rect 6906 9216 6912 9280
rect 6976 9216 6992 9280
rect 7056 9216 7072 9280
rect 7136 9216 7152 9280
rect 7216 9216 7232 9280
rect 7296 9216 7302 9280
rect 6906 9215 7302 9216
rect 10906 9280 11302 9281
rect 10906 9216 10912 9280
rect 10976 9216 10992 9280
rect 11056 9216 11072 9280
rect 11136 9216 11152 9280
rect 11216 9216 11232 9280
rect 11296 9216 11302 9280
rect 10906 9215 11302 9216
rect 14906 9280 15302 9281
rect 14906 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15072 9280
rect 15136 9216 15152 9280
rect 15216 9216 15232 9280
rect 15296 9216 15302 9280
rect 14906 9215 15302 9216
rect 18906 9280 19302 9281
rect 18906 9216 18912 9280
rect 18976 9216 18992 9280
rect 19056 9216 19072 9280
rect 19136 9216 19152 9280
rect 19216 9216 19232 9280
rect 19296 9216 19302 9280
rect 18906 9215 19302 9216
rect 22906 9280 23302 9281
rect 22906 9216 22912 9280
rect 22976 9216 22992 9280
rect 23056 9216 23072 9280
rect 23136 9216 23152 9280
rect 23216 9216 23232 9280
rect 23296 9216 23302 9280
rect 22906 9215 23302 9216
rect 3646 8736 4042 8737
rect 3646 8672 3652 8736
rect 3716 8672 3732 8736
rect 3796 8672 3812 8736
rect 3876 8672 3892 8736
rect 3956 8672 3972 8736
rect 4036 8672 4042 8736
rect 3646 8671 4042 8672
rect 7646 8736 8042 8737
rect 7646 8672 7652 8736
rect 7716 8672 7732 8736
rect 7796 8672 7812 8736
rect 7876 8672 7892 8736
rect 7956 8672 7972 8736
rect 8036 8672 8042 8736
rect 7646 8671 8042 8672
rect 11646 8736 12042 8737
rect 11646 8672 11652 8736
rect 11716 8672 11732 8736
rect 11796 8672 11812 8736
rect 11876 8672 11892 8736
rect 11956 8672 11972 8736
rect 12036 8672 12042 8736
rect 11646 8671 12042 8672
rect 15646 8736 16042 8737
rect 15646 8672 15652 8736
rect 15716 8672 15732 8736
rect 15796 8672 15812 8736
rect 15876 8672 15892 8736
rect 15956 8672 15972 8736
rect 16036 8672 16042 8736
rect 15646 8671 16042 8672
rect 19646 8736 20042 8737
rect 19646 8672 19652 8736
rect 19716 8672 19732 8736
rect 19796 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20042 8736
rect 19646 8671 20042 8672
rect 23646 8736 24042 8737
rect 23646 8672 23652 8736
rect 23716 8672 23732 8736
rect 23796 8672 23812 8736
rect 23876 8672 23892 8736
rect 23956 8672 23972 8736
rect 24036 8672 24042 8736
rect 23646 8671 24042 8672
rect 5165 8530 5231 8533
rect 10593 8530 10659 8533
rect 14549 8532 14615 8533
rect 14549 8530 14596 8532
rect 5165 8528 14596 8530
rect 14660 8530 14666 8532
rect 20713 8530 20779 8533
rect 14660 8528 20779 8530
rect 5165 8472 5170 8528
rect 5226 8472 10598 8528
rect 10654 8472 14554 8528
rect 14660 8472 20718 8528
rect 20774 8472 20779 8528
rect 5165 8470 14596 8472
rect 5165 8467 5231 8470
rect 10593 8467 10659 8470
rect 14549 8468 14596 8470
rect 14660 8470 20779 8472
rect 14660 8468 14666 8470
rect 14549 8467 14615 8468
rect 20713 8467 20779 8470
rect 2906 8192 3302 8193
rect 2906 8128 2912 8192
rect 2976 8128 2992 8192
rect 3056 8128 3072 8192
rect 3136 8128 3152 8192
rect 3216 8128 3232 8192
rect 3296 8128 3302 8192
rect 2906 8127 3302 8128
rect 6906 8192 7302 8193
rect 6906 8128 6912 8192
rect 6976 8128 6992 8192
rect 7056 8128 7072 8192
rect 7136 8128 7152 8192
rect 7216 8128 7232 8192
rect 7296 8128 7302 8192
rect 6906 8127 7302 8128
rect 10906 8192 11302 8193
rect 10906 8128 10912 8192
rect 10976 8128 10992 8192
rect 11056 8128 11072 8192
rect 11136 8128 11152 8192
rect 11216 8128 11232 8192
rect 11296 8128 11302 8192
rect 10906 8127 11302 8128
rect 14906 8192 15302 8193
rect 14906 8128 14912 8192
rect 14976 8128 14992 8192
rect 15056 8128 15072 8192
rect 15136 8128 15152 8192
rect 15216 8128 15232 8192
rect 15296 8128 15302 8192
rect 14906 8127 15302 8128
rect 18906 8192 19302 8193
rect 18906 8128 18912 8192
rect 18976 8128 18992 8192
rect 19056 8128 19072 8192
rect 19136 8128 19152 8192
rect 19216 8128 19232 8192
rect 19296 8128 19302 8192
rect 18906 8127 19302 8128
rect 22906 8192 23302 8193
rect 22906 8128 22912 8192
rect 22976 8128 22992 8192
rect 23056 8128 23072 8192
rect 23136 8128 23152 8192
rect 23216 8128 23232 8192
rect 23296 8128 23302 8192
rect 22906 8127 23302 8128
rect 18638 7924 18644 7988
rect 18708 7986 18714 7988
rect 19701 7986 19767 7989
rect 18708 7984 19767 7986
rect 18708 7928 19706 7984
rect 19762 7928 19767 7984
rect 18708 7926 19767 7928
rect 18708 7924 18714 7926
rect 19701 7923 19767 7926
rect 11237 7850 11303 7853
rect 15377 7850 15443 7853
rect 11237 7848 15443 7850
rect 11237 7792 11242 7848
rect 11298 7792 15382 7848
rect 15438 7792 15443 7848
rect 11237 7790 15443 7792
rect 11237 7787 11303 7790
rect 15377 7787 15443 7790
rect 3646 7648 4042 7649
rect 3646 7584 3652 7648
rect 3716 7584 3732 7648
rect 3796 7584 3812 7648
rect 3876 7584 3892 7648
rect 3956 7584 3972 7648
rect 4036 7584 4042 7648
rect 3646 7583 4042 7584
rect 7646 7648 8042 7649
rect 7646 7584 7652 7648
rect 7716 7584 7732 7648
rect 7796 7584 7812 7648
rect 7876 7584 7892 7648
rect 7956 7584 7972 7648
rect 8036 7584 8042 7648
rect 7646 7583 8042 7584
rect 11646 7648 12042 7649
rect 11646 7584 11652 7648
rect 11716 7584 11732 7648
rect 11796 7584 11812 7648
rect 11876 7584 11892 7648
rect 11956 7584 11972 7648
rect 12036 7584 12042 7648
rect 11646 7583 12042 7584
rect 15646 7648 16042 7649
rect 15646 7584 15652 7648
rect 15716 7584 15732 7648
rect 15796 7584 15812 7648
rect 15876 7584 15892 7648
rect 15956 7584 15972 7648
rect 16036 7584 16042 7648
rect 15646 7583 16042 7584
rect 19646 7648 20042 7649
rect 19646 7584 19652 7648
rect 19716 7584 19732 7648
rect 19796 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20042 7648
rect 19646 7583 20042 7584
rect 23646 7648 24042 7649
rect 23646 7584 23652 7648
rect 23716 7584 23732 7648
rect 23796 7584 23812 7648
rect 23876 7584 23892 7648
rect 23956 7584 23972 7648
rect 24036 7584 24042 7648
rect 23646 7583 24042 7584
rect 26509 7578 26575 7581
rect 27171 7578 27971 7608
rect 26509 7576 27971 7578
rect 26509 7520 26514 7576
rect 26570 7520 27971 7576
rect 26509 7518 27971 7520
rect 26509 7515 26575 7518
rect 27171 7488 27971 7518
rect 3601 7442 3667 7445
rect 4521 7442 4587 7445
rect 3601 7440 4587 7442
rect 3601 7384 3606 7440
rect 3662 7384 4526 7440
rect 4582 7384 4587 7440
rect 3601 7382 4587 7384
rect 3601 7379 3667 7382
rect 4521 7379 4587 7382
rect 5717 7442 5783 7445
rect 7741 7442 7807 7445
rect 8293 7442 8359 7445
rect 5717 7440 8359 7442
rect 5717 7384 5722 7440
rect 5778 7384 7746 7440
rect 7802 7384 8298 7440
rect 8354 7384 8359 7440
rect 5717 7382 8359 7384
rect 5717 7379 5783 7382
rect 7741 7379 7807 7382
rect 8293 7379 8359 7382
rect 21633 7306 21699 7309
rect 26325 7306 26391 7309
rect 21633 7304 26391 7306
rect 21633 7248 21638 7304
rect 21694 7248 26330 7304
rect 26386 7248 26391 7304
rect 21633 7246 26391 7248
rect 21633 7243 21699 7246
rect 26325 7243 26391 7246
rect 2906 7104 3302 7105
rect 2906 7040 2912 7104
rect 2976 7040 2992 7104
rect 3056 7040 3072 7104
rect 3136 7040 3152 7104
rect 3216 7040 3232 7104
rect 3296 7040 3302 7104
rect 2906 7039 3302 7040
rect 6906 7104 7302 7105
rect 6906 7040 6912 7104
rect 6976 7040 6992 7104
rect 7056 7040 7072 7104
rect 7136 7040 7152 7104
rect 7216 7040 7232 7104
rect 7296 7040 7302 7104
rect 6906 7039 7302 7040
rect 10906 7104 11302 7105
rect 10906 7040 10912 7104
rect 10976 7040 10992 7104
rect 11056 7040 11072 7104
rect 11136 7040 11152 7104
rect 11216 7040 11232 7104
rect 11296 7040 11302 7104
rect 10906 7039 11302 7040
rect 14906 7104 15302 7105
rect 14906 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15072 7104
rect 15136 7040 15152 7104
rect 15216 7040 15232 7104
rect 15296 7040 15302 7104
rect 14906 7039 15302 7040
rect 18906 7104 19302 7105
rect 18906 7040 18912 7104
rect 18976 7040 18992 7104
rect 19056 7040 19072 7104
rect 19136 7040 19152 7104
rect 19216 7040 19232 7104
rect 19296 7040 19302 7104
rect 18906 7039 19302 7040
rect 22906 7104 23302 7105
rect 22906 7040 22912 7104
rect 22976 7040 22992 7104
rect 23056 7040 23072 7104
rect 23136 7040 23152 7104
rect 23216 7040 23232 7104
rect 23296 7040 23302 7104
rect 22906 7039 23302 7040
rect 5165 7036 5231 7037
rect 5165 7034 5212 7036
rect 5120 7032 5212 7034
rect 5120 6976 5170 7032
rect 5120 6974 5212 6976
rect 5165 6972 5212 6974
rect 5276 6972 5282 7036
rect 5165 6971 5231 6972
rect 18045 6762 18111 6765
rect 18454 6762 18460 6764
rect 18045 6760 18460 6762
rect 18045 6704 18050 6760
rect 18106 6704 18460 6760
rect 18045 6702 18460 6704
rect 18045 6699 18111 6702
rect 18454 6700 18460 6702
rect 18524 6762 18530 6764
rect 20989 6762 21055 6765
rect 18524 6760 21055 6762
rect 18524 6704 20994 6760
rect 21050 6704 21055 6760
rect 18524 6702 21055 6704
rect 18524 6700 18530 6702
rect 20989 6699 21055 6702
rect 3646 6560 4042 6561
rect 3646 6496 3652 6560
rect 3716 6496 3732 6560
rect 3796 6496 3812 6560
rect 3876 6496 3892 6560
rect 3956 6496 3972 6560
rect 4036 6496 4042 6560
rect 3646 6495 4042 6496
rect 7646 6560 8042 6561
rect 7646 6496 7652 6560
rect 7716 6496 7732 6560
rect 7796 6496 7812 6560
rect 7876 6496 7892 6560
rect 7956 6496 7972 6560
rect 8036 6496 8042 6560
rect 7646 6495 8042 6496
rect 11646 6560 12042 6561
rect 11646 6496 11652 6560
rect 11716 6496 11732 6560
rect 11796 6496 11812 6560
rect 11876 6496 11892 6560
rect 11956 6496 11972 6560
rect 12036 6496 12042 6560
rect 11646 6495 12042 6496
rect 15646 6560 16042 6561
rect 15646 6496 15652 6560
rect 15716 6496 15732 6560
rect 15796 6496 15812 6560
rect 15876 6496 15892 6560
rect 15956 6496 15972 6560
rect 16036 6496 16042 6560
rect 15646 6495 16042 6496
rect 19646 6560 20042 6561
rect 19646 6496 19652 6560
rect 19716 6496 19732 6560
rect 19796 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20042 6560
rect 19646 6495 20042 6496
rect 23646 6560 24042 6561
rect 23646 6496 23652 6560
rect 23716 6496 23732 6560
rect 23796 6496 23812 6560
rect 23876 6496 23892 6560
rect 23956 6496 23972 6560
rect 24036 6496 24042 6560
rect 23646 6495 24042 6496
rect 20897 6354 20963 6357
rect 22093 6354 22159 6357
rect 20897 6352 22159 6354
rect 20897 6296 20902 6352
rect 20958 6296 22098 6352
rect 22154 6296 22159 6352
rect 20897 6294 22159 6296
rect 20897 6291 20963 6294
rect 22093 6291 22159 6294
rect 25405 6354 25471 6357
rect 25957 6354 26023 6357
rect 25405 6352 26023 6354
rect 25405 6296 25410 6352
rect 25466 6296 25962 6352
rect 26018 6296 26023 6352
rect 25405 6294 26023 6296
rect 25405 6291 25471 6294
rect 25957 6291 26023 6294
rect 2906 6016 3302 6017
rect 2906 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3072 6016
rect 3136 5952 3152 6016
rect 3216 5952 3232 6016
rect 3296 5952 3302 6016
rect 2906 5951 3302 5952
rect 6906 6016 7302 6017
rect 6906 5952 6912 6016
rect 6976 5952 6992 6016
rect 7056 5952 7072 6016
rect 7136 5952 7152 6016
rect 7216 5952 7232 6016
rect 7296 5952 7302 6016
rect 6906 5951 7302 5952
rect 10906 6016 11302 6017
rect 10906 5952 10912 6016
rect 10976 5952 10992 6016
rect 11056 5952 11072 6016
rect 11136 5952 11152 6016
rect 11216 5952 11232 6016
rect 11296 5952 11302 6016
rect 10906 5951 11302 5952
rect 14906 6016 15302 6017
rect 14906 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15072 6016
rect 15136 5952 15152 6016
rect 15216 5952 15232 6016
rect 15296 5952 15302 6016
rect 14906 5951 15302 5952
rect 18906 6016 19302 6017
rect 18906 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19302 6016
rect 18906 5951 19302 5952
rect 22906 6016 23302 6017
rect 22906 5952 22912 6016
rect 22976 5952 22992 6016
rect 23056 5952 23072 6016
rect 23136 5952 23152 6016
rect 23216 5952 23232 6016
rect 23296 5952 23302 6016
rect 22906 5951 23302 5952
rect 3646 5472 4042 5473
rect 3646 5408 3652 5472
rect 3716 5408 3732 5472
rect 3796 5408 3812 5472
rect 3876 5408 3892 5472
rect 3956 5408 3972 5472
rect 4036 5408 4042 5472
rect 3646 5407 4042 5408
rect 7646 5472 8042 5473
rect 7646 5408 7652 5472
rect 7716 5408 7732 5472
rect 7796 5408 7812 5472
rect 7876 5408 7892 5472
rect 7956 5408 7972 5472
rect 8036 5408 8042 5472
rect 7646 5407 8042 5408
rect 11646 5472 12042 5473
rect 11646 5408 11652 5472
rect 11716 5408 11732 5472
rect 11796 5408 11812 5472
rect 11876 5408 11892 5472
rect 11956 5408 11972 5472
rect 12036 5408 12042 5472
rect 11646 5407 12042 5408
rect 15646 5472 16042 5473
rect 15646 5408 15652 5472
rect 15716 5408 15732 5472
rect 15796 5408 15812 5472
rect 15876 5408 15892 5472
rect 15956 5408 15972 5472
rect 16036 5408 16042 5472
rect 15646 5407 16042 5408
rect 19646 5472 20042 5473
rect 19646 5408 19652 5472
rect 19716 5408 19732 5472
rect 19796 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20042 5472
rect 19646 5407 20042 5408
rect 23646 5472 24042 5473
rect 23646 5408 23652 5472
rect 23716 5408 23732 5472
rect 23796 5408 23812 5472
rect 23876 5408 23892 5472
rect 23956 5408 23972 5472
rect 24036 5408 24042 5472
rect 23646 5407 24042 5408
rect 2906 4928 3302 4929
rect 2906 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3072 4928
rect 3136 4864 3152 4928
rect 3216 4864 3232 4928
rect 3296 4864 3302 4928
rect 2906 4863 3302 4864
rect 6906 4928 7302 4929
rect 6906 4864 6912 4928
rect 6976 4864 6992 4928
rect 7056 4864 7072 4928
rect 7136 4864 7152 4928
rect 7216 4864 7232 4928
rect 7296 4864 7302 4928
rect 6906 4863 7302 4864
rect 10906 4928 11302 4929
rect 10906 4864 10912 4928
rect 10976 4864 10992 4928
rect 11056 4864 11072 4928
rect 11136 4864 11152 4928
rect 11216 4864 11232 4928
rect 11296 4864 11302 4928
rect 10906 4863 11302 4864
rect 14906 4928 15302 4929
rect 14906 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15072 4928
rect 15136 4864 15152 4928
rect 15216 4864 15232 4928
rect 15296 4864 15302 4928
rect 14906 4863 15302 4864
rect 18906 4928 19302 4929
rect 18906 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19302 4928
rect 18906 4863 19302 4864
rect 22906 4928 23302 4929
rect 22906 4864 22912 4928
rect 22976 4864 22992 4928
rect 23056 4864 23072 4928
rect 23136 4864 23152 4928
rect 23216 4864 23232 4928
rect 23296 4864 23302 4928
rect 22906 4863 23302 4864
rect 3646 4384 4042 4385
rect 3646 4320 3652 4384
rect 3716 4320 3732 4384
rect 3796 4320 3812 4384
rect 3876 4320 3892 4384
rect 3956 4320 3972 4384
rect 4036 4320 4042 4384
rect 3646 4319 4042 4320
rect 7646 4384 8042 4385
rect 7646 4320 7652 4384
rect 7716 4320 7732 4384
rect 7796 4320 7812 4384
rect 7876 4320 7892 4384
rect 7956 4320 7972 4384
rect 8036 4320 8042 4384
rect 7646 4319 8042 4320
rect 11646 4384 12042 4385
rect 11646 4320 11652 4384
rect 11716 4320 11732 4384
rect 11796 4320 11812 4384
rect 11876 4320 11892 4384
rect 11956 4320 11972 4384
rect 12036 4320 12042 4384
rect 11646 4319 12042 4320
rect 15646 4384 16042 4385
rect 15646 4320 15652 4384
rect 15716 4320 15732 4384
rect 15796 4320 15812 4384
rect 15876 4320 15892 4384
rect 15956 4320 15972 4384
rect 16036 4320 16042 4384
rect 15646 4319 16042 4320
rect 19646 4384 20042 4385
rect 19646 4320 19652 4384
rect 19716 4320 19732 4384
rect 19796 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20042 4384
rect 19646 4319 20042 4320
rect 23646 4384 24042 4385
rect 23646 4320 23652 4384
rect 23716 4320 23732 4384
rect 23796 4320 23812 4384
rect 23876 4320 23892 4384
rect 23956 4320 23972 4384
rect 24036 4320 24042 4384
rect 23646 4319 24042 4320
rect 2906 3840 3302 3841
rect 2906 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3072 3840
rect 3136 3776 3152 3840
rect 3216 3776 3232 3840
rect 3296 3776 3302 3840
rect 2906 3775 3302 3776
rect 6906 3840 7302 3841
rect 6906 3776 6912 3840
rect 6976 3776 6992 3840
rect 7056 3776 7072 3840
rect 7136 3776 7152 3840
rect 7216 3776 7232 3840
rect 7296 3776 7302 3840
rect 6906 3775 7302 3776
rect 10906 3840 11302 3841
rect 10906 3776 10912 3840
rect 10976 3776 10992 3840
rect 11056 3776 11072 3840
rect 11136 3776 11152 3840
rect 11216 3776 11232 3840
rect 11296 3776 11302 3840
rect 10906 3775 11302 3776
rect 14906 3840 15302 3841
rect 14906 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15072 3840
rect 15136 3776 15152 3840
rect 15216 3776 15232 3840
rect 15296 3776 15302 3840
rect 14906 3775 15302 3776
rect 18906 3840 19302 3841
rect 18906 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19302 3840
rect 18906 3775 19302 3776
rect 22906 3840 23302 3841
rect 22906 3776 22912 3840
rect 22976 3776 22992 3840
rect 23056 3776 23072 3840
rect 23136 3776 23152 3840
rect 23216 3776 23232 3840
rect 23296 3776 23302 3840
rect 22906 3775 23302 3776
rect 3646 3296 4042 3297
rect 3646 3232 3652 3296
rect 3716 3232 3732 3296
rect 3796 3232 3812 3296
rect 3876 3232 3892 3296
rect 3956 3232 3972 3296
rect 4036 3232 4042 3296
rect 3646 3231 4042 3232
rect 7646 3296 8042 3297
rect 7646 3232 7652 3296
rect 7716 3232 7732 3296
rect 7796 3232 7812 3296
rect 7876 3232 7892 3296
rect 7956 3232 7972 3296
rect 8036 3232 8042 3296
rect 7646 3231 8042 3232
rect 11646 3296 12042 3297
rect 11646 3232 11652 3296
rect 11716 3232 11732 3296
rect 11796 3232 11812 3296
rect 11876 3232 11892 3296
rect 11956 3232 11972 3296
rect 12036 3232 12042 3296
rect 11646 3231 12042 3232
rect 15646 3296 16042 3297
rect 15646 3232 15652 3296
rect 15716 3232 15732 3296
rect 15796 3232 15812 3296
rect 15876 3232 15892 3296
rect 15956 3232 15972 3296
rect 16036 3232 16042 3296
rect 15646 3231 16042 3232
rect 19646 3296 20042 3297
rect 19646 3232 19652 3296
rect 19716 3232 19732 3296
rect 19796 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20042 3296
rect 19646 3231 20042 3232
rect 23646 3296 24042 3297
rect 23646 3232 23652 3296
rect 23716 3232 23732 3296
rect 23796 3232 23812 3296
rect 23876 3232 23892 3296
rect 23956 3232 23972 3296
rect 24036 3232 24042 3296
rect 23646 3231 24042 3232
rect 2906 2752 3302 2753
rect 2906 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3072 2752
rect 3136 2688 3152 2752
rect 3216 2688 3232 2752
rect 3296 2688 3302 2752
rect 2906 2687 3302 2688
rect 6906 2752 7302 2753
rect 6906 2688 6912 2752
rect 6976 2688 6992 2752
rect 7056 2688 7072 2752
rect 7136 2688 7152 2752
rect 7216 2688 7232 2752
rect 7296 2688 7302 2752
rect 6906 2687 7302 2688
rect 10906 2752 11302 2753
rect 10906 2688 10912 2752
rect 10976 2688 10992 2752
rect 11056 2688 11072 2752
rect 11136 2688 11152 2752
rect 11216 2688 11232 2752
rect 11296 2688 11302 2752
rect 10906 2687 11302 2688
rect 14906 2752 15302 2753
rect 14906 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15072 2752
rect 15136 2688 15152 2752
rect 15216 2688 15232 2752
rect 15296 2688 15302 2752
rect 14906 2687 15302 2688
rect 18906 2752 19302 2753
rect 18906 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19302 2752
rect 18906 2687 19302 2688
rect 22906 2752 23302 2753
rect 22906 2688 22912 2752
rect 22976 2688 22992 2752
rect 23056 2688 23072 2752
rect 23136 2688 23152 2752
rect 23216 2688 23232 2752
rect 23296 2688 23302 2752
rect 22906 2687 23302 2688
rect 3646 2208 4042 2209
rect 3646 2144 3652 2208
rect 3716 2144 3732 2208
rect 3796 2144 3812 2208
rect 3876 2144 3892 2208
rect 3956 2144 3972 2208
rect 4036 2144 4042 2208
rect 3646 2143 4042 2144
rect 7646 2208 8042 2209
rect 7646 2144 7652 2208
rect 7716 2144 7732 2208
rect 7796 2144 7812 2208
rect 7876 2144 7892 2208
rect 7956 2144 7972 2208
rect 8036 2144 8042 2208
rect 7646 2143 8042 2144
rect 11646 2208 12042 2209
rect 11646 2144 11652 2208
rect 11716 2144 11732 2208
rect 11796 2144 11812 2208
rect 11876 2144 11892 2208
rect 11956 2144 11972 2208
rect 12036 2144 12042 2208
rect 11646 2143 12042 2144
rect 15646 2208 16042 2209
rect 15646 2144 15652 2208
rect 15716 2144 15732 2208
rect 15796 2144 15812 2208
rect 15876 2144 15892 2208
rect 15956 2144 15972 2208
rect 16036 2144 16042 2208
rect 15646 2143 16042 2144
rect 19646 2208 20042 2209
rect 19646 2144 19652 2208
rect 19716 2144 19732 2208
rect 19796 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20042 2208
rect 19646 2143 20042 2144
rect 23646 2208 24042 2209
rect 23646 2144 23652 2208
rect 23716 2144 23732 2208
rect 23796 2144 23812 2208
rect 23876 2144 23892 2208
rect 23956 2144 23972 2208
rect 24036 2144 24042 2208
rect 23646 2143 24042 2144
<< via3 >>
rect 2912 27772 2976 27776
rect 2912 27716 2916 27772
rect 2916 27716 2972 27772
rect 2972 27716 2976 27772
rect 2912 27712 2976 27716
rect 2992 27772 3056 27776
rect 2992 27716 2996 27772
rect 2996 27716 3052 27772
rect 3052 27716 3056 27772
rect 2992 27712 3056 27716
rect 3072 27772 3136 27776
rect 3072 27716 3076 27772
rect 3076 27716 3132 27772
rect 3132 27716 3136 27772
rect 3072 27712 3136 27716
rect 3152 27772 3216 27776
rect 3152 27716 3156 27772
rect 3156 27716 3212 27772
rect 3212 27716 3216 27772
rect 3152 27712 3216 27716
rect 3232 27772 3296 27776
rect 3232 27716 3236 27772
rect 3236 27716 3292 27772
rect 3292 27716 3296 27772
rect 3232 27712 3296 27716
rect 6912 27772 6976 27776
rect 6912 27716 6916 27772
rect 6916 27716 6972 27772
rect 6972 27716 6976 27772
rect 6912 27712 6976 27716
rect 6992 27772 7056 27776
rect 6992 27716 6996 27772
rect 6996 27716 7052 27772
rect 7052 27716 7056 27772
rect 6992 27712 7056 27716
rect 7072 27772 7136 27776
rect 7072 27716 7076 27772
rect 7076 27716 7132 27772
rect 7132 27716 7136 27772
rect 7072 27712 7136 27716
rect 7152 27772 7216 27776
rect 7152 27716 7156 27772
rect 7156 27716 7212 27772
rect 7212 27716 7216 27772
rect 7152 27712 7216 27716
rect 7232 27772 7296 27776
rect 7232 27716 7236 27772
rect 7236 27716 7292 27772
rect 7292 27716 7296 27772
rect 7232 27712 7296 27716
rect 10912 27772 10976 27776
rect 10912 27716 10916 27772
rect 10916 27716 10972 27772
rect 10972 27716 10976 27772
rect 10912 27712 10976 27716
rect 10992 27772 11056 27776
rect 10992 27716 10996 27772
rect 10996 27716 11052 27772
rect 11052 27716 11056 27772
rect 10992 27712 11056 27716
rect 11072 27772 11136 27776
rect 11072 27716 11076 27772
rect 11076 27716 11132 27772
rect 11132 27716 11136 27772
rect 11072 27712 11136 27716
rect 11152 27772 11216 27776
rect 11152 27716 11156 27772
rect 11156 27716 11212 27772
rect 11212 27716 11216 27772
rect 11152 27712 11216 27716
rect 11232 27772 11296 27776
rect 11232 27716 11236 27772
rect 11236 27716 11292 27772
rect 11292 27716 11296 27772
rect 11232 27712 11296 27716
rect 14912 27772 14976 27776
rect 14912 27716 14916 27772
rect 14916 27716 14972 27772
rect 14972 27716 14976 27772
rect 14912 27712 14976 27716
rect 14992 27772 15056 27776
rect 14992 27716 14996 27772
rect 14996 27716 15052 27772
rect 15052 27716 15056 27772
rect 14992 27712 15056 27716
rect 15072 27772 15136 27776
rect 15072 27716 15076 27772
rect 15076 27716 15132 27772
rect 15132 27716 15136 27772
rect 15072 27712 15136 27716
rect 15152 27772 15216 27776
rect 15152 27716 15156 27772
rect 15156 27716 15212 27772
rect 15212 27716 15216 27772
rect 15152 27712 15216 27716
rect 15232 27772 15296 27776
rect 15232 27716 15236 27772
rect 15236 27716 15292 27772
rect 15292 27716 15296 27772
rect 15232 27712 15296 27716
rect 18912 27772 18976 27776
rect 18912 27716 18916 27772
rect 18916 27716 18972 27772
rect 18972 27716 18976 27772
rect 18912 27712 18976 27716
rect 18992 27772 19056 27776
rect 18992 27716 18996 27772
rect 18996 27716 19052 27772
rect 19052 27716 19056 27772
rect 18992 27712 19056 27716
rect 19072 27772 19136 27776
rect 19072 27716 19076 27772
rect 19076 27716 19132 27772
rect 19132 27716 19136 27772
rect 19072 27712 19136 27716
rect 19152 27772 19216 27776
rect 19152 27716 19156 27772
rect 19156 27716 19212 27772
rect 19212 27716 19216 27772
rect 19152 27712 19216 27716
rect 19232 27772 19296 27776
rect 19232 27716 19236 27772
rect 19236 27716 19292 27772
rect 19292 27716 19296 27772
rect 19232 27712 19296 27716
rect 22912 27772 22976 27776
rect 22912 27716 22916 27772
rect 22916 27716 22972 27772
rect 22972 27716 22976 27772
rect 22912 27712 22976 27716
rect 22992 27772 23056 27776
rect 22992 27716 22996 27772
rect 22996 27716 23052 27772
rect 23052 27716 23056 27772
rect 22992 27712 23056 27716
rect 23072 27772 23136 27776
rect 23072 27716 23076 27772
rect 23076 27716 23132 27772
rect 23132 27716 23136 27772
rect 23072 27712 23136 27716
rect 23152 27772 23216 27776
rect 23152 27716 23156 27772
rect 23156 27716 23212 27772
rect 23212 27716 23216 27772
rect 23152 27712 23216 27716
rect 23232 27772 23296 27776
rect 23232 27716 23236 27772
rect 23236 27716 23292 27772
rect 23292 27716 23296 27772
rect 23232 27712 23296 27716
rect 3652 27228 3716 27232
rect 3652 27172 3656 27228
rect 3656 27172 3712 27228
rect 3712 27172 3716 27228
rect 3652 27168 3716 27172
rect 3732 27228 3796 27232
rect 3732 27172 3736 27228
rect 3736 27172 3792 27228
rect 3792 27172 3796 27228
rect 3732 27168 3796 27172
rect 3812 27228 3876 27232
rect 3812 27172 3816 27228
rect 3816 27172 3872 27228
rect 3872 27172 3876 27228
rect 3812 27168 3876 27172
rect 3892 27228 3956 27232
rect 3892 27172 3896 27228
rect 3896 27172 3952 27228
rect 3952 27172 3956 27228
rect 3892 27168 3956 27172
rect 3972 27228 4036 27232
rect 3972 27172 3976 27228
rect 3976 27172 4032 27228
rect 4032 27172 4036 27228
rect 3972 27168 4036 27172
rect 7652 27228 7716 27232
rect 7652 27172 7656 27228
rect 7656 27172 7712 27228
rect 7712 27172 7716 27228
rect 7652 27168 7716 27172
rect 7732 27228 7796 27232
rect 7732 27172 7736 27228
rect 7736 27172 7792 27228
rect 7792 27172 7796 27228
rect 7732 27168 7796 27172
rect 7812 27228 7876 27232
rect 7812 27172 7816 27228
rect 7816 27172 7872 27228
rect 7872 27172 7876 27228
rect 7812 27168 7876 27172
rect 7892 27228 7956 27232
rect 7892 27172 7896 27228
rect 7896 27172 7952 27228
rect 7952 27172 7956 27228
rect 7892 27168 7956 27172
rect 7972 27228 8036 27232
rect 7972 27172 7976 27228
rect 7976 27172 8032 27228
rect 8032 27172 8036 27228
rect 7972 27168 8036 27172
rect 11652 27228 11716 27232
rect 11652 27172 11656 27228
rect 11656 27172 11712 27228
rect 11712 27172 11716 27228
rect 11652 27168 11716 27172
rect 11732 27228 11796 27232
rect 11732 27172 11736 27228
rect 11736 27172 11792 27228
rect 11792 27172 11796 27228
rect 11732 27168 11796 27172
rect 11812 27228 11876 27232
rect 11812 27172 11816 27228
rect 11816 27172 11872 27228
rect 11872 27172 11876 27228
rect 11812 27168 11876 27172
rect 11892 27228 11956 27232
rect 11892 27172 11896 27228
rect 11896 27172 11952 27228
rect 11952 27172 11956 27228
rect 11892 27168 11956 27172
rect 11972 27228 12036 27232
rect 11972 27172 11976 27228
rect 11976 27172 12032 27228
rect 12032 27172 12036 27228
rect 11972 27168 12036 27172
rect 15652 27228 15716 27232
rect 15652 27172 15656 27228
rect 15656 27172 15712 27228
rect 15712 27172 15716 27228
rect 15652 27168 15716 27172
rect 15732 27228 15796 27232
rect 15732 27172 15736 27228
rect 15736 27172 15792 27228
rect 15792 27172 15796 27228
rect 15732 27168 15796 27172
rect 15812 27228 15876 27232
rect 15812 27172 15816 27228
rect 15816 27172 15872 27228
rect 15872 27172 15876 27228
rect 15812 27168 15876 27172
rect 15892 27228 15956 27232
rect 15892 27172 15896 27228
rect 15896 27172 15952 27228
rect 15952 27172 15956 27228
rect 15892 27168 15956 27172
rect 15972 27228 16036 27232
rect 15972 27172 15976 27228
rect 15976 27172 16032 27228
rect 16032 27172 16036 27228
rect 15972 27168 16036 27172
rect 19652 27228 19716 27232
rect 19652 27172 19656 27228
rect 19656 27172 19712 27228
rect 19712 27172 19716 27228
rect 19652 27168 19716 27172
rect 19732 27228 19796 27232
rect 19732 27172 19736 27228
rect 19736 27172 19792 27228
rect 19792 27172 19796 27228
rect 19732 27168 19796 27172
rect 19812 27228 19876 27232
rect 19812 27172 19816 27228
rect 19816 27172 19872 27228
rect 19872 27172 19876 27228
rect 19812 27168 19876 27172
rect 19892 27228 19956 27232
rect 19892 27172 19896 27228
rect 19896 27172 19952 27228
rect 19952 27172 19956 27228
rect 19892 27168 19956 27172
rect 19972 27228 20036 27232
rect 19972 27172 19976 27228
rect 19976 27172 20032 27228
rect 20032 27172 20036 27228
rect 19972 27168 20036 27172
rect 23652 27228 23716 27232
rect 23652 27172 23656 27228
rect 23656 27172 23712 27228
rect 23712 27172 23716 27228
rect 23652 27168 23716 27172
rect 23732 27228 23796 27232
rect 23732 27172 23736 27228
rect 23736 27172 23792 27228
rect 23792 27172 23796 27228
rect 23732 27168 23796 27172
rect 23812 27228 23876 27232
rect 23812 27172 23816 27228
rect 23816 27172 23872 27228
rect 23872 27172 23876 27228
rect 23812 27168 23876 27172
rect 23892 27228 23956 27232
rect 23892 27172 23896 27228
rect 23896 27172 23952 27228
rect 23952 27172 23956 27228
rect 23892 27168 23956 27172
rect 23972 27228 24036 27232
rect 23972 27172 23976 27228
rect 23976 27172 24032 27228
rect 24032 27172 24036 27228
rect 23972 27168 24036 27172
rect 10180 26828 10244 26892
rect 2912 26684 2976 26688
rect 2912 26628 2916 26684
rect 2916 26628 2972 26684
rect 2972 26628 2976 26684
rect 2912 26624 2976 26628
rect 2992 26684 3056 26688
rect 2992 26628 2996 26684
rect 2996 26628 3052 26684
rect 3052 26628 3056 26684
rect 2992 26624 3056 26628
rect 3072 26684 3136 26688
rect 3072 26628 3076 26684
rect 3076 26628 3132 26684
rect 3132 26628 3136 26684
rect 3072 26624 3136 26628
rect 3152 26684 3216 26688
rect 3152 26628 3156 26684
rect 3156 26628 3212 26684
rect 3212 26628 3216 26684
rect 3152 26624 3216 26628
rect 3232 26684 3296 26688
rect 3232 26628 3236 26684
rect 3236 26628 3292 26684
rect 3292 26628 3296 26684
rect 3232 26624 3296 26628
rect 6912 26684 6976 26688
rect 6912 26628 6916 26684
rect 6916 26628 6972 26684
rect 6972 26628 6976 26684
rect 6912 26624 6976 26628
rect 6992 26684 7056 26688
rect 6992 26628 6996 26684
rect 6996 26628 7052 26684
rect 7052 26628 7056 26684
rect 6992 26624 7056 26628
rect 7072 26684 7136 26688
rect 7072 26628 7076 26684
rect 7076 26628 7132 26684
rect 7132 26628 7136 26684
rect 7072 26624 7136 26628
rect 7152 26684 7216 26688
rect 7152 26628 7156 26684
rect 7156 26628 7212 26684
rect 7212 26628 7216 26684
rect 7152 26624 7216 26628
rect 7232 26684 7296 26688
rect 7232 26628 7236 26684
rect 7236 26628 7292 26684
rect 7292 26628 7296 26684
rect 7232 26624 7296 26628
rect 10912 26684 10976 26688
rect 10912 26628 10916 26684
rect 10916 26628 10972 26684
rect 10972 26628 10976 26684
rect 10912 26624 10976 26628
rect 10992 26684 11056 26688
rect 10992 26628 10996 26684
rect 10996 26628 11052 26684
rect 11052 26628 11056 26684
rect 10992 26624 11056 26628
rect 11072 26684 11136 26688
rect 11072 26628 11076 26684
rect 11076 26628 11132 26684
rect 11132 26628 11136 26684
rect 11072 26624 11136 26628
rect 11152 26684 11216 26688
rect 11152 26628 11156 26684
rect 11156 26628 11212 26684
rect 11212 26628 11216 26684
rect 11152 26624 11216 26628
rect 11232 26684 11296 26688
rect 11232 26628 11236 26684
rect 11236 26628 11292 26684
rect 11292 26628 11296 26684
rect 11232 26624 11296 26628
rect 14912 26684 14976 26688
rect 14912 26628 14916 26684
rect 14916 26628 14972 26684
rect 14972 26628 14976 26684
rect 14912 26624 14976 26628
rect 14992 26684 15056 26688
rect 14992 26628 14996 26684
rect 14996 26628 15052 26684
rect 15052 26628 15056 26684
rect 14992 26624 15056 26628
rect 15072 26684 15136 26688
rect 15072 26628 15076 26684
rect 15076 26628 15132 26684
rect 15132 26628 15136 26684
rect 15072 26624 15136 26628
rect 15152 26684 15216 26688
rect 15152 26628 15156 26684
rect 15156 26628 15212 26684
rect 15212 26628 15216 26684
rect 15152 26624 15216 26628
rect 15232 26684 15296 26688
rect 15232 26628 15236 26684
rect 15236 26628 15292 26684
rect 15292 26628 15296 26684
rect 15232 26624 15296 26628
rect 18912 26684 18976 26688
rect 18912 26628 18916 26684
rect 18916 26628 18972 26684
rect 18972 26628 18976 26684
rect 18912 26624 18976 26628
rect 18992 26684 19056 26688
rect 18992 26628 18996 26684
rect 18996 26628 19052 26684
rect 19052 26628 19056 26684
rect 18992 26624 19056 26628
rect 19072 26684 19136 26688
rect 19072 26628 19076 26684
rect 19076 26628 19132 26684
rect 19132 26628 19136 26684
rect 19072 26624 19136 26628
rect 19152 26684 19216 26688
rect 19152 26628 19156 26684
rect 19156 26628 19212 26684
rect 19212 26628 19216 26684
rect 19152 26624 19216 26628
rect 19232 26684 19296 26688
rect 19232 26628 19236 26684
rect 19236 26628 19292 26684
rect 19292 26628 19296 26684
rect 19232 26624 19296 26628
rect 22912 26684 22976 26688
rect 22912 26628 22916 26684
rect 22916 26628 22972 26684
rect 22972 26628 22976 26684
rect 22912 26624 22976 26628
rect 22992 26684 23056 26688
rect 22992 26628 22996 26684
rect 22996 26628 23052 26684
rect 23052 26628 23056 26684
rect 22992 26624 23056 26628
rect 23072 26684 23136 26688
rect 23072 26628 23076 26684
rect 23076 26628 23132 26684
rect 23132 26628 23136 26684
rect 23072 26624 23136 26628
rect 23152 26684 23216 26688
rect 23152 26628 23156 26684
rect 23156 26628 23212 26684
rect 23212 26628 23216 26684
rect 23152 26624 23216 26628
rect 23232 26684 23296 26688
rect 23232 26628 23236 26684
rect 23236 26628 23292 26684
rect 23292 26628 23296 26684
rect 23232 26624 23296 26628
rect 3652 26140 3716 26144
rect 3652 26084 3656 26140
rect 3656 26084 3712 26140
rect 3712 26084 3716 26140
rect 3652 26080 3716 26084
rect 3732 26140 3796 26144
rect 3732 26084 3736 26140
rect 3736 26084 3792 26140
rect 3792 26084 3796 26140
rect 3732 26080 3796 26084
rect 3812 26140 3876 26144
rect 3812 26084 3816 26140
rect 3816 26084 3872 26140
rect 3872 26084 3876 26140
rect 3812 26080 3876 26084
rect 3892 26140 3956 26144
rect 3892 26084 3896 26140
rect 3896 26084 3952 26140
rect 3952 26084 3956 26140
rect 3892 26080 3956 26084
rect 3972 26140 4036 26144
rect 3972 26084 3976 26140
rect 3976 26084 4032 26140
rect 4032 26084 4036 26140
rect 3972 26080 4036 26084
rect 7652 26140 7716 26144
rect 7652 26084 7656 26140
rect 7656 26084 7712 26140
rect 7712 26084 7716 26140
rect 7652 26080 7716 26084
rect 7732 26140 7796 26144
rect 7732 26084 7736 26140
rect 7736 26084 7792 26140
rect 7792 26084 7796 26140
rect 7732 26080 7796 26084
rect 7812 26140 7876 26144
rect 7812 26084 7816 26140
rect 7816 26084 7872 26140
rect 7872 26084 7876 26140
rect 7812 26080 7876 26084
rect 7892 26140 7956 26144
rect 7892 26084 7896 26140
rect 7896 26084 7952 26140
rect 7952 26084 7956 26140
rect 7892 26080 7956 26084
rect 7972 26140 8036 26144
rect 7972 26084 7976 26140
rect 7976 26084 8032 26140
rect 8032 26084 8036 26140
rect 7972 26080 8036 26084
rect 11652 26140 11716 26144
rect 11652 26084 11656 26140
rect 11656 26084 11712 26140
rect 11712 26084 11716 26140
rect 11652 26080 11716 26084
rect 11732 26140 11796 26144
rect 11732 26084 11736 26140
rect 11736 26084 11792 26140
rect 11792 26084 11796 26140
rect 11732 26080 11796 26084
rect 11812 26140 11876 26144
rect 11812 26084 11816 26140
rect 11816 26084 11872 26140
rect 11872 26084 11876 26140
rect 11812 26080 11876 26084
rect 11892 26140 11956 26144
rect 11892 26084 11896 26140
rect 11896 26084 11952 26140
rect 11952 26084 11956 26140
rect 11892 26080 11956 26084
rect 11972 26140 12036 26144
rect 11972 26084 11976 26140
rect 11976 26084 12032 26140
rect 12032 26084 12036 26140
rect 11972 26080 12036 26084
rect 15652 26140 15716 26144
rect 15652 26084 15656 26140
rect 15656 26084 15712 26140
rect 15712 26084 15716 26140
rect 15652 26080 15716 26084
rect 15732 26140 15796 26144
rect 15732 26084 15736 26140
rect 15736 26084 15792 26140
rect 15792 26084 15796 26140
rect 15732 26080 15796 26084
rect 15812 26140 15876 26144
rect 15812 26084 15816 26140
rect 15816 26084 15872 26140
rect 15872 26084 15876 26140
rect 15812 26080 15876 26084
rect 15892 26140 15956 26144
rect 15892 26084 15896 26140
rect 15896 26084 15952 26140
rect 15952 26084 15956 26140
rect 15892 26080 15956 26084
rect 15972 26140 16036 26144
rect 15972 26084 15976 26140
rect 15976 26084 16032 26140
rect 16032 26084 16036 26140
rect 15972 26080 16036 26084
rect 19652 26140 19716 26144
rect 19652 26084 19656 26140
rect 19656 26084 19712 26140
rect 19712 26084 19716 26140
rect 19652 26080 19716 26084
rect 19732 26140 19796 26144
rect 19732 26084 19736 26140
rect 19736 26084 19792 26140
rect 19792 26084 19796 26140
rect 19732 26080 19796 26084
rect 19812 26140 19876 26144
rect 19812 26084 19816 26140
rect 19816 26084 19872 26140
rect 19872 26084 19876 26140
rect 19812 26080 19876 26084
rect 19892 26140 19956 26144
rect 19892 26084 19896 26140
rect 19896 26084 19952 26140
rect 19952 26084 19956 26140
rect 19892 26080 19956 26084
rect 19972 26140 20036 26144
rect 19972 26084 19976 26140
rect 19976 26084 20032 26140
rect 20032 26084 20036 26140
rect 19972 26080 20036 26084
rect 23652 26140 23716 26144
rect 23652 26084 23656 26140
rect 23656 26084 23712 26140
rect 23712 26084 23716 26140
rect 23652 26080 23716 26084
rect 23732 26140 23796 26144
rect 23732 26084 23736 26140
rect 23736 26084 23792 26140
rect 23792 26084 23796 26140
rect 23732 26080 23796 26084
rect 23812 26140 23876 26144
rect 23812 26084 23816 26140
rect 23816 26084 23872 26140
rect 23872 26084 23876 26140
rect 23812 26080 23876 26084
rect 23892 26140 23956 26144
rect 23892 26084 23896 26140
rect 23896 26084 23952 26140
rect 23952 26084 23956 26140
rect 23892 26080 23956 26084
rect 23972 26140 24036 26144
rect 23972 26084 23976 26140
rect 23976 26084 24032 26140
rect 24032 26084 24036 26140
rect 23972 26080 24036 26084
rect 2912 25596 2976 25600
rect 2912 25540 2916 25596
rect 2916 25540 2972 25596
rect 2972 25540 2976 25596
rect 2912 25536 2976 25540
rect 2992 25596 3056 25600
rect 2992 25540 2996 25596
rect 2996 25540 3052 25596
rect 3052 25540 3056 25596
rect 2992 25536 3056 25540
rect 3072 25596 3136 25600
rect 3072 25540 3076 25596
rect 3076 25540 3132 25596
rect 3132 25540 3136 25596
rect 3072 25536 3136 25540
rect 3152 25596 3216 25600
rect 3152 25540 3156 25596
rect 3156 25540 3212 25596
rect 3212 25540 3216 25596
rect 3152 25536 3216 25540
rect 3232 25596 3296 25600
rect 3232 25540 3236 25596
rect 3236 25540 3292 25596
rect 3292 25540 3296 25596
rect 3232 25536 3296 25540
rect 6912 25596 6976 25600
rect 6912 25540 6916 25596
rect 6916 25540 6972 25596
rect 6972 25540 6976 25596
rect 6912 25536 6976 25540
rect 6992 25596 7056 25600
rect 6992 25540 6996 25596
rect 6996 25540 7052 25596
rect 7052 25540 7056 25596
rect 6992 25536 7056 25540
rect 7072 25596 7136 25600
rect 7072 25540 7076 25596
rect 7076 25540 7132 25596
rect 7132 25540 7136 25596
rect 7072 25536 7136 25540
rect 7152 25596 7216 25600
rect 7152 25540 7156 25596
rect 7156 25540 7212 25596
rect 7212 25540 7216 25596
rect 7152 25536 7216 25540
rect 7232 25596 7296 25600
rect 7232 25540 7236 25596
rect 7236 25540 7292 25596
rect 7292 25540 7296 25596
rect 7232 25536 7296 25540
rect 10912 25596 10976 25600
rect 10912 25540 10916 25596
rect 10916 25540 10972 25596
rect 10972 25540 10976 25596
rect 10912 25536 10976 25540
rect 10992 25596 11056 25600
rect 10992 25540 10996 25596
rect 10996 25540 11052 25596
rect 11052 25540 11056 25596
rect 10992 25536 11056 25540
rect 11072 25596 11136 25600
rect 11072 25540 11076 25596
rect 11076 25540 11132 25596
rect 11132 25540 11136 25596
rect 11072 25536 11136 25540
rect 11152 25596 11216 25600
rect 11152 25540 11156 25596
rect 11156 25540 11212 25596
rect 11212 25540 11216 25596
rect 11152 25536 11216 25540
rect 11232 25596 11296 25600
rect 11232 25540 11236 25596
rect 11236 25540 11292 25596
rect 11292 25540 11296 25596
rect 11232 25536 11296 25540
rect 14912 25596 14976 25600
rect 14912 25540 14916 25596
rect 14916 25540 14972 25596
rect 14972 25540 14976 25596
rect 14912 25536 14976 25540
rect 14992 25596 15056 25600
rect 14992 25540 14996 25596
rect 14996 25540 15052 25596
rect 15052 25540 15056 25596
rect 14992 25536 15056 25540
rect 15072 25596 15136 25600
rect 15072 25540 15076 25596
rect 15076 25540 15132 25596
rect 15132 25540 15136 25596
rect 15072 25536 15136 25540
rect 15152 25596 15216 25600
rect 15152 25540 15156 25596
rect 15156 25540 15212 25596
rect 15212 25540 15216 25596
rect 15152 25536 15216 25540
rect 15232 25596 15296 25600
rect 15232 25540 15236 25596
rect 15236 25540 15292 25596
rect 15292 25540 15296 25596
rect 15232 25536 15296 25540
rect 18912 25596 18976 25600
rect 18912 25540 18916 25596
rect 18916 25540 18972 25596
rect 18972 25540 18976 25596
rect 18912 25536 18976 25540
rect 18992 25596 19056 25600
rect 18992 25540 18996 25596
rect 18996 25540 19052 25596
rect 19052 25540 19056 25596
rect 18992 25536 19056 25540
rect 19072 25596 19136 25600
rect 19072 25540 19076 25596
rect 19076 25540 19132 25596
rect 19132 25540 19136 25596
rect 19072 25536 19136 25540
rect 19152 25596 19216 25600
rect 19152 25540 19156 25596
rect 19156 25540 19212 25596
rect 19212 25540 19216 25596
rect 19152 25536 19216 25540
rect 19232 25596 19296 25600
rect 19232 25540 19236 25596
rect 19236 25540 19292 25596
rect 19292 25540 19296 25596
rect 19232 25536 19296 25540
rect 22912 25596 22976 25600
rect 22912 25540 22916 25596
rect 22916 25540 22972 25596
rect 22972 25540 22976 25596
rect 22912 25536 22976 25540
rect 22992 25596 23056 25600
rect 22992 25540 22996 25596
rect 22996 25540 23052 25596
rect 23052 25540 23056 25596
rect 22992 25536 23056 25540
rect 23072 25596 23136 25600
rect 23072 25540 23076 25596
rect 23076 25540 23132 25596
rect 23132 25540 23136 25596
rect 23072 25536 23136 25540
rect 23152 25596 23216 25600
rect 23152 25540 23156 25596
rect 23156 25540 23212 25596
rect 23212 25540 23216 25596
rect 23152 25536 23216 25540
rect 23232 25596 23296 25600
rect 23232 25540 23236 25596
rect 23236 25540 23292 25596
rect 23292 25540 23296 25596
rect 23232 25536 23296 25540
rect 3652 25052 3716 25056
rect 3652 24996 3656 25052
rect 3656 24996 3712 25052
rect 3712 24996 3716 25052
rect 3652 24992 3716 24996
rect 3732 25052 3796 25056
rect 3732 24996 3736 25052
rect 3736 24996 3792 25052
rect 3792 24996 3796 25052
rect 3732 24992 3796 24996
rect 3812 25052 3876 25056
rect 3812 24996 3816 25052
rect 3816 24996 3872 25052
rect 3872 24996 3876 25052
rect 3812 24992 3876 24996
rect 3892 25052 3956 25056
rect 3892 24996 3896 25052
rect 3896 24996 3952 25052
rect 3952 24996 3956 25052
rect 3892 24992 3956 24996
rect 3972 25052 4036 25056
rect 3972 24996 3976 25052
rect 3976 24996 4032 25052
rect 4032 24996 4036 25052
rect 3972 24992 4036 24996
rect 7652 25052 7716 25056
rect 7652 24996 7656 25052
rect 7656 24996 7712 25052
rect 7712 24996 7716 25052
rect 7652 24992 7716 24996
rect 7732 25052 7796 25056
rect 7732 24996 7736 25052
rect 7736 24996 7792 25052
rect 7792 24996 7796 25052
rect 7732 24992 7796 24996
rect 7812 25052 7876 25056
rect 7812 24996 7816 25052
rect 7816 24996 7872 25052
rect 7872 24996 7876 25052
rect 7812 24992 7876 24996
rect 7892 25052 7956 25056
rect 7892 24996 7896 25052
rect 7896 24996 7952 25052
rect 7952 24996 7956 25052
rect 7892 24992 7956 24996
rect 7972 25052 8036 25056
rect 7972 24996 7976 25052
rect 7976 24996 8032 25052
rect 8032 24996 8036 25052
rect 7972 24992 8036 24996
rect 11652 25052 11716 25056
rect 11652 24996 11656 25052
rect 11656 24996 11712 25052
rect 11712 24996 11716 25052
rect 11652 24992 11716 24996
rect 11732 25052 11796 25056
rect 11732 24996 11736 25052
rect 11736 24996 11792 25052
rect 11792 24996 11796 25052
rect 11732 24992 11796 24996
rect 11812 25052 11876 25056
rect 11812 24996 11816 25052
rect 11816 24996 11872 25052
rect 11872 24996 11876 25052
rect 11812 24992 11876 24996
rect 11892 25052 11956 25056
rect 11892 24996 11896 25052
rect 11896 24996 11952 25052
rect 11952 24996 11956 25052
rect 11892 24992 11956 24996
rect 11972 25052 12036 25056
rect 11972 24996 11976 25052
rect 11976 24996 12032 25052
rect 12032 24996 12036 25052
rect 11972 24992 12036 24996
rect 15652 25052 15716 25056
rect 15652 24996 15656 25052
rect 15656 24996 15712 25052
rect 15712 24996 15716 25052
rect 15652 24992 15716 24996
rect 15732 25052 15796 25056
rect 15732 24996 15736 25052
rect 15736 24996 15792 25052
rect 15792 24996 15796 25052
rect 15732 24992 15796 24996
rect 15812 25052 15876 25056
rect 15812 24996 15816 25052
rect 15816 24996 15872 25052
rect 15872 24996 15876 25052
rect 15812 24992 15876 24996
rect 15892 25052 15956 25056
rect 15892 24996 15896 25052
rect 15896 24996 15952 25052
rect 15952 24996 15956 25052
rect 15892 24992 15956 24996
rect 15972 25052 16036 25056
rect 15972 24996 15976 25052
rect 15976 24996 16032 25052
rect 16032 24996 16036 25052
rect 15972 24992 16036 24996
rect 19652 25052 19716 25056
rect 19652 24996 19656 25052
rect 19656 24996 19712 25052
rect 19712 24996 19716 25052
rect 19652 24992 19716 24996
rect 19732 25052 19796 25056
rect 19732 24996 19736 25052
rect 19736 24996 19792 25052
rect 19792 24996 19796 25052
rect 19732 24992 19796 24996
rect 19812 25052 19876 25056
rect 19812 24996 19816 25052
rect 19816 24996 19872 25052
rect 19872 24996 19876 25052
rect 19812 24992 19876 24996
rect 19892 25052 19956 25056
rect 19892 24996 19896 25052
rect 19896 24996 19952 25052
rect 19952 24996 19956 25052
rect 19892 24992 19956 24996
rect 19972 25052 20036 25056
rect 19972 24996 19976 25052
rect 19976 24996 20032 25052
rect 20032 24996 20036 25052
rect 19972 24992 20036 24996
rect 23652 25052 23716 25056
rect 23652 24996 23656 25052
rect 23656 24996 23712 25052
rect 23712 24996 23716 25052
rect 23652 24992 23716 24996
rect 23732 25052 23796 25056
rect 23732 24996 23736 25052
rect 23736 24996 23792 25052
rect 23792 24996 23796 25052
rect 23732 24992 23796 24996
rect 23812 25052 23876 25056
rect 23812 24996 23816 25052
rect 23816 24996 23872 25052
rect 23872 24996 23876 25052
rect 23812 24992 23876 24996
rect 23892 25052 23956 25056
rect 23892 24996 23896 25052
rect 23896 24996 23952 25052
rect 23952 24996 23956 25052
rect 23892 24992 23956 24996
rect 23972 25052 24036 25056
rect 23972 24996 23976 25052
rect 23976 24996 24032 25052
rect 24032 24996 24036 25052
rect 23972 24992 24036 24996
rect 17540 24924 17604 24988
rect 24348 24924 24412 24988
rect 2912 24508 2976 24512
rect 2912 24452 2916 24508
rect 2916 24452 2972 24508
rect 2972 24452 2976 24508
rect 2912 24448 2976 24452
rect 2992 24508 3056 24512
rect 2992 24452 2996 24508
rect 2996 24452 3052 24508
rect 3052 24452 3056 24508
rect 2992 24448 3056 24452
rect 3072 24508 3136 24512
rect 3072 24452 3076 24508
rect 3076 24452 3132 24508
rect 3132 24452 3136 24508
rect 3072 24448 3136 24452
rect 3152 24508 3216 24512
rect 3152 24452 3156 24508
rect 3156 24452 3212 24508
rect 3212 24452 3216 24508
rect 3152 24448 3216 24452
rect 3232 24508 3296 24512
rect 3232 24452 3236 24508
rect 3236 24452 3292 24508
rect 3292 24452 3296 24508
rect 3232 24448 3296 24452
rect 6912 24508 6976 24512
rect 6912 24452 6916 24508
rect 6916 24452 6972 24508
rect 6972 24452 6976 24508
rect 6912 24448 6976 24452
rect 6992 24508 7056 24512
rect 6992 24452 6996 24508
rect 6996 24452 7052 24508
rect 7052 24452 7056 24508
rect 6992 24448 7056 24452
rect 7072 24508 7136 24512
rect 7072 24452 7076 24508
rect 7076 24452 7132 24508
rect 7132 24452 7136 24508
rect 7072 24448 7136 24452
rect 7152 24508 7216 24512
rect 7152 24452 7156 24508
rect 7156 24452 7212 24508
rect 7212 24452 7216 24508
rect 7152 24448 7216 24452
rect 7232 24508 7296 24512
rect 7232 24452 7236 24508
rect 7236 24452 7292 24508
rect 7292 24452 7296 24508
rect 7232 24448 7296 24452
rect 10912 24508 10976 24512
rect 10912 24452 10916 24508
rect 10916 24452 10972 24508
rect 10972 24452 10976 24508
rect 10912 24448 10976 24452
rect 10992 24508 11056 24512
rect 10992 24452 10996 24508
rect 10996 24452 11052 24508
rect 11052 24452 11056 24508
rect 10992 24448 11056 24452
rect 11072 24508 11136 24512
rect 11072 24452 11076 24508
rect 11076 24452 11132 24508
rect 11132 24452 11136 24508
rect 11072 24448 11136 24452
rect 11152 24508 11216 24512
rect 11152 24452 11156 24508
rect 11156 24452 11212 24508
rect 11212 24452 11216 24508
rect 11152 24448 11216 24452
rect 11232 24508 11296 24512
rect 11232 24452 11236 24508
rect 11236 24452 11292 24508
rect 11292 24452 11296 24508
rect 11232 24448 11296 24452
rect 14912 24508 14976 24512
rect 14912 24452 14916 24508
rect 14916 24452 14972 24508
rect 14972 24452 14976 24508
rect 14912 24448 14976 24452
rect 14992 24508 15056 24512
rect 14992 24452 14996 24508
rect 14996 24452 15052 24508
rect 15052 24452 15056 24508
rect 14992 24448 15056 24452
rect 15072 24508 15136 24512
rect 15072 24452 15076 24508
rect 15076 24452 15132 24508
rect 15132 24452 15136 24508
rect 15072 24448 15136 24452
rect 15152 24508 15216 24512
rect 15152 24452 15156 24508
rect 15156 24452 15212 24508
rect 15212 24452 15216 24508
rect 15152 24448 15216 24452
rect 15232 24508 15296 24512
rect 15232 24452 15236 24508
rect 15236 24452 15292 24508
rect 15292 24452 15296 24508
rect 15232 24448 15296 24452
rect 18912 24508 18976 24512
rect 18912 24452 18916 24508
rect 18916 24452 18972 24508
rect 18972 24452 18976 24508
rect 18912 24448 18976 24452
rect 18992 24508 19056 24512
rect 18992 24452 18996 24508
rect 18996 24452 19052 24508
rect 19052 24452 19056 24508
rect 18992 24448 19056 24452
rect 19072 24508 19136 24512
rect 19072 24452 19076 24508
rect 19076 24452 19132 24508
rect 19132 24452 19136 24508
rect 19072 24448 19136 24452
rect 19152 24508 19216 24512
rect 19152 24452 19156 24508
rect 19156 24452 19212 24508
rect 19212 24452 19216 24508
rect 19152 24448 19216 24452
rect 19232 24508 19296 24512
rect 19232 24452 19236 24508
rect 19236 24452 19292 24508
rect 19292 24452 19296 24508
rect 19232 24448 19296 24452
rect 22912 24508 22976 24512
rect 22912 24452 22916 24508
rect 22916 24452 22972 24508
rect 22972 24452 22976 24508
rect 22912 24448 22976 24452
rect 22992 24508 23056 24512
rect 22992 24452 22996 24508
rect 22996 24452 23052 24508
rect 23052 24452 23056 24508
rect 22992 24448 23056 24452
rect 23072 24508 23136 24512
rect 23072 24452 23076 24508
rect 23076 24452 23132 24508
rect 23132 24452 23136 24508
rect 23072 24448 23136 24452
rect 23152 24508 23216 24512
rect 23152 24452 23156 24508
rect 23156 24452 23212 24508
rect 23212 24452 23216 24508
rect 23152 24448 23216 24452
rect 23232 24508 23296 24512
rect 23232 24452 23236 24508
rect 23236 24452 23292 24508
rect 23292 24452 23296 24508
rect 23232 24448 23296 24452
rect 3652 23964 3716 23968
rect 3652 23908 3656 23964
rect 3656 23908 3712 23964
rect 3712 23908 3716 23964
rect 3652 23904 3716 23908
rect 3732 23964 3796 23968
rect 3732 23908 3736 23964
rect 3736 23908 3792 23964
rect 3792 23908 3796 23964
rect 3732 23904 3796 23908
rect 3812 23964 3876 23968
rect 3812 23908 3816 23964
rect 3816 23908 3872 23964
rect 3872 23908 3876 23964
rect 3812 23904 3876 23908
rect 3892 23964 3956 23968
rect 3892 23908 3896 23964
rect 3896 23908 3952 23964
rect 3952 23908 3956 23964
rect 3892 23904 3956 23908
rect 3972 23964 4036 23968
rect 3972 23908 3976 23964
rect 3976 23908 4032 23964
rect 4032 23908 4036 23964
rect 3972 23904 4036 23908
rect 7652 23964 7716 23968
rect 7652 23908 7656 23964
rect 7656 23908 7712 23964
rect 7712 23908 7716 23964
rect 7652 23904 7716 23908
rect 7732 23964 7796 23968
rect 7732 23908 7736 23964
rect 7736 23908 7792 23964
rect 7792 23908 7796 23964
rect 7732 23904 7796 23908
rect 7812 23964 7876 23968
rect 7812 23908 7816 23964
rect 7816 23908 7872 23964
rect 7872 23908 7876 23964
rect 7812 23904 7876 23908
rect 7892 23964 7956 23968
rect 7892 23908 7896 23964
rect 7896 23908 7952 23964
rect 7952 23908 7956 23964
rect 7892 23904 7956 23908
rect 7972 23964 8036 23968
rect 7972 23908 7976 23964
rect 7976 23908 8032 23964
rect 8032 23908 8036 23964
rect 7972 23904 8036 23908
rect 11652 23964 11716 23968
rect 11652 23908 11656 23964
rect 11656 23908 11712 23964
rect 11712 23908 11716 23964
rect 11652 23904 11716 23908
rect 11732 23964 11796 23968
rect 11732 23908 11736 23964
rect 11736 23908 11792 23964
rect 11792 23908 11796 23964
rect 11732 23904 11796 23908
rect 11812 23964 11876 23968
rect 11812 23908 11816 23964
rect 11816 23908 11872 23964
rect 11872 23908 11876 23964
rect 11812 23904 11876 23908
rect 11892 23964 11956 23968
rect 11892 23908 11896 23964
rect 11896 23908 11952 23964
rect 11952 23908 11956 23964
rect 11892 23904 11956 23908
rect 11972 23964 12036 23968
rect 11972 23908 11976 23964
rect 11976 23908 12032 23964
rect 12032 23908 12036 23964
rect 11972 23904 12036 23908
rect 15652 23964 15716 23968
rect 15652 23908 15656 23964
rect 15656 23908 15712 23964
rect 15712 23908 15716 23964
rect 15652 23904 15716 23908
rect 15732 23964 15796 23968
rect 15732 23908 15736 23964
rect 15736 23908 15792 23964
rect 15792 23908 15796 23964
rect 15732 23904 15796 23908
rect 15812 23964 15876 23968
rect 15812 23908 15816 23964
rect 15816 23908 15872 23964
rect 15872 23908 15876 23964
rect 15812 23904 15876 23908
rect 15892 23964 15956 23968
rect 15892 23908 15896 23964
rect 15896 23908 15952 23964
rect 15952 23908 15956 23964
rect 15892 23904 15956 23908
rect 15972 23964 16036 23968
rect 15972 23908 15976 23964
rect 15976 23908 16032 23964
rect 16032 23908 16036 23964
rect 15972 23904 16036 23908
rect 19652 23964 19716 23968
rect 19652 23908 19656 23964
rect 19656 23908 19712 23964
rect 19712 23908 19716 23964
rect 19652 23904 19716 23908
rect 19732 23964 19796 23968
rect 19732 23908 19736 23964
rect 19736 23908 19792 23964
rect 19792 23908 19796 23964
rect 19732 23904 19796 23908
rect 19812 23964 19876 23968
rect 19812 23908 19816 23964
rect 19816 23908 19872 23964
rect 19872 23908 19876 23964
rect 19812 23904 19876 23908
rect 19892 23964 19956 23968
rect 19892 23908 19896 23964
rect 19896 23908 19952 23964
rect 19952 23908 19956 23964
rect 19892 23904 19956 23908
rect 19972 23964 20036 23968
rect 19972 23908 19976 23964
rect 19976 23908 20032 23964
rect 20032 23908 20036 23964
rect 19972 23904 20036 23908
rect 23652 23964 23716 23968
rect 23652 23908 23656 23964
rect 23656 23908 23712 23964
rect 23712 23908 23716 23964
rect 23652 23904 23716 23908
rect 23732 23964 23796 23968
rect 23732 23908 23736 23964
rect 23736 23908 23792 23964
rect 23792 23908 23796 23964
rect 23732 23904 23796 23908
rect 23812 23964 23876 23968
rect 23812 23908 23816 23964
rect 23816 23908 23872 23964
rect 23872 23908 23876 23964
rect 23812 23904 23876 23908
rect 23892 23964 23956 23968
rect 23892 23908 23896 23964
rect 23896 23908 23952 23964
rect 23952 23908 23956 23964
rect 23892 23904 23956 23908
rect 23972 23964 24036 23968
rect 23972 23908 23976 23964
rect 23976 23908 24032 23964
rect 24032 23908 24036 23964
rect 23972 23904 24036 23908
rect 2912 23420 2976 23424
rect 2912 23364 2916 23420
rect 2916 23364 2972 23420
rect 2972 23364 2976 23420
rect 2912 23360 2976 23364
rect 2992 23420 3056 23424
rect 2992 23364 2996 23420
rect 2996 23364 3052 23420
rect 3052 23364 3056 23420
rect 2992 23360 3056 23364
rect 3072 23420 3136 23424
rect 3072 23364 3076 23420
rect 3076 23364 3132 23420
rect 3132 23364 3136 23420
rect 3072 23360 3136 23364
rect 3152 23420 3216 23424
rect 3152 23364 3156 23420
rect 3156 23364 3212 23420
rect 3212 23364 3216 23420
rect 3152 23360 3216 23364
rect 3232 23420 3296 23424
rect 3232 23364 3236 23420
rect 3236 23364 3292 23420
rect 3292 23364 3296 23420
rect 3232 23360 3296 23364
rect 6912 23420 6976 23424
rect 6912 23364 6916 23420
rect 6916 23364 6972 23420
rect 6972 23364 6976 23420
rect 6912 23360 6976 23364
rect 6992 23420 7056 23424
rect 6992 23364 6996 23420
rect 6996 23364 7052 23420
rect 7052 23364 7056 23420
rect 6992 23360 7056 23364
rect 7072 23420 7136 23424
rect 7072 23364 7076 23420
rect 7076 23364 7132 23420
rect 7132 23364 7136 23420
rect 7072 23360 7136 23364
rect 7152 23420 7216 23424
rect 7152 23364 7156 23420
rect 7156 23364 7212 23420
rect 7212 23364 7216 23420
rect 7152 23360 7216 23364
rect 7232 23420 7296 23424
rect 7232 23364 7236 23420
rect 7236 23364 7292 23420
rect 7292 23364 7296 23420
rect 7232 23360 7296 23364
rect 10912 23420 10976 23424
rect 10912 23364 10916 23420
rect 10916 23364 10972 23420
rect 10972 23364 10976 23420
rect 10912 23360 10976 23364
rect 10992 23420 11056 23424
rect 10992 23364 10996 23420
rect 10996 23364 11052 23420
rect 11052 23364 11056 23420
rect 10992 23360 11056 23364
rect 11072 23420 11136 23424
rect 11072 23364 11076 23420
rect 11076 23364 11132 23420
rect 11132 23364 11136 23420
rect 11072 23360 11136 23364
rect 11152 23420 11216 23424
rect 11152 23364 11156 23420
rect 11156 23364 11212 23420
rect 11212 23364 11216 23420
rect 11152 23360 11216 23364
rect 11232 23420 11296 23424
rect 11232 23364 11236 23420
rect 11236 23364 11292 23420
rect 11292 23364 11296 23420
rect 11232 23360 11296 23364
rect 14912 23420 14976 23424
rect 14912 23364 14916 23420
rect 14916 23364 14972 23420
rect 14972 23364 14976 23420
rect 14912 23360 14976 23364
rect 14992 23420 15056 23424
rect 14992 23364 14996 23420
rect 14996 23364 15052 23420
rect 15052 23364 15056 23420
rect 14992 23360 15056 23364
rect 15072 23420 15136 23424
rect 15072 23364 15076 23420
rect 15076 23364 15132 23420
rect 15132 23364 15136 23420
rect 15072 23360 15136 23364
rect 15152 23420 15216 23424
rect 15152 23364 15156 23420
rect 15156 23364 15212 23420
rect 15212 23364 15216 23420
rect 15152 23360 15216 23364
rect 15232 23420 15296 23424
rect 15232 23364 15236 23420
rect 15236 23364 15292 23420
rect 15292 23364 15296 23420
rect 15232 23360 15296 23364
rect 18912 23420 18976 23424
rect 18912 23364 18916 23420
rect 18916 23364 18972 23420
rect 18972 23364 18976 23420
rect 18912 23360 18976 23364
rect 18992 23420 19056 23424
rect 18992 23364 18996 23420
rect 18996 23364 19052 23420
rect 19052 23364 19056 23420
rect 18992 23360 19056 23364
rect 19072 23420 19136 23424
rect 19072 23364 19076 23420
rect 19076 23364 19132 23420
rect 19132 23364 19136 23420
rect 19072 23360 19136 23364
rect 19152 23420 19216 23424
rect 19152 23364 19156 23420
rect 19156 23364 19212 23420
rect 19212 23364 19216 23420
rect 19152 23360 19216 23364
rect 19232 23420 19296 23424
rect 19232 23364 19236 23420
rect 19236 23364 19292 23420
rect 19292 23364 19296 23420
rect 19232 23360 19296 23364
rect 22912 23420 22976 23424
rect 22912 23364 22916 23420
rect 22916 23364 22972 23420
rect 22972 23364 22976 23420
rect 22912 23360 22976 23364
rect 22992 23420 23056 23424
rect 22992 23364 22996 23420
rect 22996 23364 23052 23420
rect 23052 23364 23056 23420
rect 22992 23360 23056 23364
rect 23072 23420 23136 23424
rect 23072 23364 23076 23420
rect 23076 23364 23132 23420
rect 23132 23364 23136 23420
rect 23072 23360 23136 23364
rect 23152 23420 23216 23424
rect 23152 23364 23156 23420
rect 23156 23364 23212 23420
rect 23212 23364 23216 23420
rect 23152 23360 23216 23364
rect 23232 23420 23296 23424
rect 23232 23364 23236 23420
rect 23236 23364 23292 23420
rect 23292 23364 23296 23420
rect 23232 23360 23296 23364
rect 3652 22876 3716 22880
rect 3652 22820 3656 22876
rect 3656 22820 3712 22876
rect 3712 22820 3716 22876
rect 3652 22816 3716 22820
rect 3732 22876 3796 22880
rect 3732 22820 3736 22876
rect 3736 22820 3792 22876
rect 3792 22820 3796 22876
rect 3732 22816 3796 22820
rect 3812 22876 3876 22880
rect 3812 22820 3816 22876
rect 3816 22820 3872 22876
rect 3872 22820 3876 22876
rect 3812 22816 3876 22820
rect 3892 22876 3956 22880
rect 3892 22820 3896 22876
rect 3896 22820 3952 22876
rect 3952 22820 3956 22876
rect 3892 22816 3956 22820
rect 3972 22876 4036 22880
rect 3972 22820 3976 22876
rect 3976 22820 4032 22876
rect 4032 22820 4036 22876
rect 3972 22816 4036 22820
rect 7652 22876 7716 22880
rect 7652 22820 7656 22876
rect 7656 22820 7712 22876
rect 7712 22820 7716 22876
rect 7652 22816 7716 22820
rect 7732 22876 7796 22880
rect 7732 22820 7736 22876
rect 7736 22820 7792 22876
rect 7792 22820 7796 22876
rect 7732 22816 7796 22820
rect 7812 22876 7876 22880
rect 7812 22820 7816 22876
rect 7816 22820 7872 22876
rect 7872 22820 7876 22876
rect 7812 22816 7876 22820
rect 7892 22876 7956 22880
rect 7892 22820 7896 22876
rect 7896 22820 7952 22876
rect 7952 22820 7956 22876
rect 7892 22816 7956 22820
rect 7972 22876 8036 22880
rect 7972 22820 7976 22876
rect 7976 22820 8032 22876
rect 8032 22820 8036 22876
rect 7972 22816 8036 22820
rect 11652 22876 11716 22880
rect 11652 22820 11656 22876
rect 11656 22820 11712 22876
rect 11712 22820 11716 22876
rect 11652 22816 11716 22820
rect 11732 22876 11796 22880
rect 11732 22820 11736 22876
rect 11736 22820 11792 22876
rect 11792 22820 11796 22876
rect 11732 22816 11796 22820
rect 11812 22876 11876 22880
rect 11812 22820 11816 22876
rect 11816 22820 11872 22876
rect 11872 22820 11876 22876
rect 11812 22816 11876 22820
rect 11892 22876 11956 22880
rect 11892 22820 11896 22876
rect 11896 22820 11952 22876
rect 11952 22820 11956 22876
rect 11892 22816 11956 22820
rect 11972 22876 12036 22880
rect 11972 22820 11976 22876
rect 11976 22820 12032 22876
rect 12032 22820 12036 22876
rect 11972 22816 12036 22820
rect 15652 22876 15716 22880
rect 15652 22820 15656 22876
rect 15656 22820 15712 22876
rect 15712 22820 15716 22876
rect 15652 22816 15716 22820
rect 15732 22876 15796 22880
rect 15732 22820 15736 22876
rect 15736 22820 15792 22876
rect 15792 22820 15796 22876
rect 15732 22816 15796 22820
rect 15812 22876 15876 22880
rect 15812 22820 15816 22876
rect 15816 22820 15872 22876
rect 15872 22820 15876 22876
rect 15812 22816 15876 22820
rect 15892 22876 15956 22880
rect 15892 22820 15896 22876
rect 15896 22820 15952 22876
rect 15952 22820 15956 22876
rect 15892 22816 15956 22820
rect 15972 22876 16036 22880
rect 15972 22820 15976 22876
rect 15976 22820 16032 22876
rect 16032 22820 16036 22876
rect 15972 22816 16036 22820
rect 19652 22876 19716 22880
rect 19652 22820 19656 22876
rect 19656 22820 19712 22876
rect 19712 22820 19716 22876
rect 19652 22816 19716 22820
rect 19732 22876 19796 22880
rect 19732 22820 19736 22876
rect 19736 22820 19792 22876
rect 19792 22820 19796 22876
rect 19732 22816 19796 22820
rect 19812 22876 19876 22880
rect 19812 22820 19816 22876
rect 19816 22820 19872 22876
rect 19872 22820 19876 22876
rect 19812 22816 19876 22820
rect 19892 22876 19956 22880
rect 19892 22820 19896 22876
rect 19896 22820 19952 22876
rect 19952 22820 19956 22876
rect 19892 22816 19956 22820
rect 19972 22876 20036 22880
rect 19972 22820 19976 22876
rect 19976 22820 20032 22876
rect 20032 22820 20036 22876
rect 19972 22816 20036 22820
rect 23652 22876 23716 22880
rect 23652 22820 23656 22876
rect 23656 22820 23712 22876
rect 23712 22820 23716 22876
rect 23652 22816 23716 22820
rect 23732 22876 23796 22880
rect 23732 22820 23736 22876
rect 23736 22820 23792 22876
rect 23792 22820 23796 22876
rect 23732 22816 23796 22820
rect 23812 22876 23876 22880
rect 23812 22820 23816 22876
rect 23816 22820 23872 22876
rect 23872 22820 23876 22876
rect 23812 22816 23876 22820
rect 23892 22876 23956 22880
rect 23892 22820 23896 22876
rect 23896 22820 23952 22876
rect 23952 22820 23956 22876
rect 23892 22816 23956 22820
rect 23972 22876 24036 22880
rect 23972 22820 23976 22876
rect 23976 22820 24032 22876
rect 24032 22820 24036 22876
rect 23972 22816 24036 22820
rect 17356 22476 17420 22540
rect 2912 22332 2976 22336
rect 2912 22276 2916 22332
rect 2916 22276 2972 22332
rect 2972 22276 2976 22332
rect 2912 22272 2976 22276
rect 2992 22332 3056 22336
rect 2992 22276 2996 22332
rect 2996 22276 3052 22332
rect 3052 22276 3056 22332
rect 2992 22272 3056 22276
rect 3072 22332 3136 22336
rect 3072 22276 3076 22332
rect 3076 22276 3132 22332
rect 3132 22276 3136 22332
rect 3072 22272 3136 22276
rect 3152 22332 3216 22336
rect 3152 22276 3156 22332
rect 3156 22276 3212 22332
rect 3212 22276 3216 22332
rect 3152 22272 3216 22276
rect 3232 22332 3296 22336
rect 3232 22276 3236 22332
rect 3236 22276 3292 22332
rect 3292 22276 3296 22332
rect 3232 22272 3296 22276
rect 6912 22332 6976 22336
rect 6912 22276 6916 22332
rect 6916 22276 6972 22332
rect 6972 22276 6976 22332
rect 6912 22272 6976 22276
rect 6992 22332 7056 22336
rect 6992 22276 6996 22332
rect 6996 22276 7052 22332
rect 7052 22276 7056 22332
rect 6992 22272 7056 22276
rect 7072 22332 7136 22336
rect 7072 22276 7076 22332
rect 7076 22276 7132 22332
rect 7132 22276 7136 22332
rect 7072 22272 7136 22276
rect 7152 22332 7216 22336
rect 7152 22276 7156 22332
rect 7156 22276 7212 22332
rect 7212 22276 7216 22332
rect 7152 22272 7216 22276
rect 7232 22332 7296 22336
rect 7232 22276 7236 22332
rect 7236 22276 7292 22332
rect 7292 22276 7296 22332
rect 7232 22272 7296 22276
rect 10912 22332 10976 22336
rect 10912 22276 10916 22332
rect 10916 22276 10972 22332
rect 10972 22276 10976 22332
rect 10912 22272 10976 22276
rect 10992 22332 11056 22336
rect 10992 22276 10996 22332
rect 10996 22276 11052 22332
rect 11052 22276 11056 22332
rect 10992 22272 11056 22276
rect 11072 22332 11136 22336
rect 11072 22276 11076 22332
rect 11076 22276 11132 22332
rect 11132 22276 11136 22332
rect 11072 22272 11136 22276
rect 11152 22332 11216 22336
rect 11152 22276 11156 22332
rect 11156 22276 11212 22332
rect 11212 22276 11216 22332
rect 11152 22272 11216 22276
rect 11232 22332 11296 22336
rect 11232 22276 11236 22332
rect 11236 22276 11292 22332
rect 11292 22276 11296 22332
rect 11232 22272 11296 22276
rect 14912 22332 14976 22336
rect 14912 22276 14916 22332
rect 14916 22276 14972 22332
rect 14972 22276 14976 22332
rect 14912 22272 14976 22276
rect 14992 22332 15056 22336
rect 14992 22276 14996 22332
rect 14996 22276 15052 22332
rect 15052 22276 15056 22332
rect 14992 22272 15056 22276
rect 15072 22332 15136 22336
rect 15072 22276 15076 22332
rect 15076 22276 15132 22332
rect 15132 22276 15136 22332
rect 15072 22272 15136 22276
rect 15152 22332 15216 22336
rect 15152 22276 15156 22332
rect 15156 22276 15212 22332
rect 15212 22276 15216 22332
rect 15152 22272 15216 22276
rect 15232 22332 15296 22336
rect 15232 22276 15236 22332
rect 15236 22276 15292 22332
rect 15292 22276 15296 22332
rect 15232 22272 15296 22276
rect 18912 22332 18976 22336
rect 18912 22276 18916 22332
rect 18916 22276 18972 22332
rect 18972 22276 18976 22332
rect 18912 22272 18976 22276
rect 18992 22332 19056 22336
rect 18992 22276 18996 22332
rect 18996 22276 19052 22332
rect 19052 22276 19056 22332
rect 18992 22272 19056 22276
rect 19072 22332 19136 22336
rect 19072 22276 19076 22332
rect 19076 22276 19132 22332
rect 19132 22276 19136 22332
rect 19072 22272 19136 22276
rect 19152 22332 19216 22336
rect 19152 22276 19156 22332
rect 19156 22276 19212 22332
rect 19212 22276 19216 22332
rect 19152 22272 19216 22276
rect 19232 22332 19296 22336
rect 19232 22276 19236 22332
rect 19236 22276 19292 22332
rect 19292 22276 19296 22332
rect 19232 22272 19296 22276
rect 22912 22332 22976 22336
rect 22912 22276 22916 22332
rect 22916 22276 22972 22332
rect 22972 22276 22976 22332
rect 22912 22272 22976 22276
rect 22992 22332 23056 22336
rect 22992 22276 22996 22332
rect 22996 22276 23052 22332
rect 23052 22276 23056 22332
rect 22992 22272 23056 22276
rect 23072 22332 23136 22336
rect 23072 22276 23076 22332
rect 23076 22276 23132 22332
rect 23132 22276 23136 22332
rect 23072 22272 23136 22276
rect 23152 22332 23216 22336
rect 23152 22276 23156 22332
rect 23156 22276 23212 22332
rect 23212 22276 23216 22332
rect 23152 22272 23216 22276
rect 23232 22332 23296 22336
rect 23232 22276 23236 22332
rect 23236 22276 23292 22332
rect 23292 22276 23296 22332
rect 23232 22272 23296 22276
rect 5396 22128 5460 22132
rect 5396 22072 5410 22128
rect 5410 22072 5460 22128
rect 5396 22068 5460 22072
rect 24348 21932 24412 21996
rect 3652 21788 3716 21792
rect 3652 21732 3656 21788
rect 3656 21732 3712 21788
rect 3712 21732 3716 21788
rect 3652 21728 3716 21732
rect 3732 21788 3796 21792
rect 3732 21732 3736 21788
rect 3736 21732 3792 21788
rect 3792 21732 3796 21788
rect 3732 21728 3796 21732
rect 3812 21788 3876 21792
rect 3812 21732 3816 21788
rect 3816 21732 3872 21788
rect 3872 21732 3876 21788
rect 3812 21728 3876 21732
rect 3892 21788 3956 21792
rect 3892 21732 3896 21788
rect 3896 21732 3952 21788
rect 3952 21732 3956 21788
rect 3892 21728 3956 21732
rect 3972 21788 4036 21792
rect 3972 21732 3976 21788
rect 3976 21732 4032 21788
rect 4032 21732 4036 21788
rect 3972 21728 4036 21732
rect 7652 21788 7716 21792
rect 7652 21732 7656 21788
rect 7656 21732 7712 21788
rect 7712 21732 7716 21788
rect 7652 21728 7716 21732
rect 7732 21788 7796 21792
rect 7732 21732 7736 21788
rect 7736 21732 7792 21788
rect 7792 21732 7796 21788
rect 7732 21728 7796 21732
rect 7812 21788 7876 21792
rect 7812 21732 7816 21788
rect 7816 21732 7872 21788
rect 7872 21732 7876 21788
rect 7812 21728 7876 21732
rect 7892 21788 7956 21792
rect 7892 21732 7896 21788
rect 7896 21732 7952 21788
rect 7952 21732 7956 21788
rect 7892 21728 7956 21732
rect 7972 21788 8036 21792
rect 7972 21732 7976 21788
rect 7976 21732 8032 21788
rect 8032 21732 8036 21788
rect 7972 21728 8036 21732
rect 11652 21788 11716 21792
rect 11652 21732 11656 21788
rect 11656 21732 11712 21788
rect 11712 21732 11716 21788
rect 11652 21728 11716 21732
rect 11732 21788 11796 21792
rect 11732 21732 11736 21788
rect 11736 21732 11792 21788
rect 11792 21732 11796 21788
rect 11732 21728 11796 21732
rect 11812 21788 11876 21792
rect 11812 21732 11816 21788
rect 11816 21732 11872 21788
rect 11872 21732 11876 21788
rect 11812 21728 11876 21732
rect 11892 21788 11956 21792
rect 11892 21732 11896 21788
rect 11896 21732 11952 21788
rect 11952 21732 11956 21788
rect 11892 21728 11956 21732
rect 11972 21788 12036 21792
rect 11972 21732 11976 21788
rect 11976 21732 12032 21788
rect 12032 21732 12036 21788
rect 11972 21728 12036 21732
rect 15652 21788 15716 21792
rect 15652 21732 15656 21788
rect 15656 21732 15712 21788
rect 15712 21732 15716 21788
rect 15652 21728 15716 21732
rect 15732 21788 15796 21792
rect 15732 21732 15736 21788
rect 15736 21732 15792 21788
rect 15792 21732 15796 21788
rect 15732 21728 15796 21732
rect 15812 21788 15876 21792
rect 15812 21732 15816 21788
rect 15816 21732 15872 21788
rect 15872 21732 15876 21788
rect 15812 21728 15876 21732
rect 15892 21788 15956 21792
rect 15892 21732 15896 21788
rect 15896 21732 15952 21788
rect 15952 21732 15956 21788
rect 15892 21728 15956 21732
rect 15972 21788 16036 21792
rect 15972 21732 15976 21788
rect 15976 21732 16032 21788
rect 16032 21732 16036 21788
rect 15972 21728 16036 21732
rect 19652 21788 19716 21792
rect 19652 21732 19656 21788
rect 19656 21732 19712 21788
rect 19712 21732 19716 21788
rect 19652 21728 19716 21732
rect 19732 21788 19796 21792
rect 19732 21732 19736 21788
rect 19736 21732 19792 21788
rect 19792 21732 19796 21788
rect 19732 21728 19796 21732
rect 19812 21788 19876 21792
rect 19812 21732 19816 21788
rect 19816 21732 19872 21788
rect 19872 21732 19876 21788
rect 19812 21728 19876 21732
rect 19892 21788 19956 21792
rect 19892 21732 19896 21788
rect 19896 21732 19952 21788
rect 19952 21732 19956 21788
rect 19892 21728 19956 21732
rect 19972 21788 20036 21792
rect 19972 21732 19976 21788
rect 19976 21732 20032 21788
rect 20032 21732 20036 21788
rect 19972 21728 20036 21732
rect 23652 21788 23716 21792
rect 23652 21732 23656 21788
rect 23656 21732 23712 21788
rect 23712 21732 23716 21788
rect 23652 21728 23716 21732
rect 23732 21788 23796 21792
rect 23732 21732 23736 21788
rect 23736 21732 23792 21788
rect 23792 21732 23796 21788
rect 23732 21728 23796 21732
rect 23812 21788 23876 21792
rect 23812 21732 23816 21788
rect 23816 21732 23872 21788
rect 23872 21732 23876 21788
rect 23812 21728 23876 21732
rect 23892 21788 23956 21792
rect 23892 21732 23896 21788
rect 23896 21732 23952 21788
rect 23952 21732 23956 21788
rect 23892 21728 23956 21732
rect 23972 21788 24036 21792
rect 23972 21732 23976 21788
rect 23976 21732 24032 21788
rect 24032 21732 24036 21788
rect 23972 21728 24036 21732
rect 2912 21244 2976 21248
rect 2912 21188 2916 21244
rect 2916 21188 2972 21244
rect 2972 21188 2976 21244
rect 2912 21184 2976 21188
rect 2992 21244 3056 21248
rect 2992 21188 2996 21244
rect 2996 21188 3052 21244
rect 3052 21188 3056 21244
rect 2992 21184 3056 21188
rect 3072 21244 3136 21248
rect 3072 21188 3076 21244
rect 3076 21188 3132 21244
rect 3132 21188 3136 21244
rect 3072 21184 3136 21188
rect 3152 21244 3216 21248
rect 3152 21188 3156 21244
rect 3156 21188 3212 21244
rect 3212 21188 3216 21244
rect 3152 21184 3216 21188
rect 3232 21244 3296 21248
rect 3232 21188 3236 21244
rect 3236 21188 3292 21244
rect 3292 21188 3296 21244
rect 3232 21184 3296 21188
rect 6912 21244 6976 21248
rect 6912 21188 6916 21244
rect 6916 21188 6972 21244
rect 6972 21188 6976 21244
rect 6912 21184 6976 21188
rect 6992 21244 7056 21248
rect 6992 21188 6996 21244
rect 6996 21188 7052 21244
rect 7052 21188 7056 21244
rect 6992 21184 7056 21188
rect 7072 21244 7136 21248
rect 7072 21188 7076 21244
rect 7076 21188 7132 21244
rect 7132 21188 7136 21244
rect 7072 21184 7136 21188
rect 7152 21244 7216 21248
rect 7152 21188 7156 21244
rect 7156 21188 7212 21244
rect 7212 21188 7216 21244
rect 7152 21184 7216 21188
rect 7232 21244 7296 21248
rect 7232 21188 7236 21244
rect 7236 21188 7292 21244
rect 7292 21188 7296 21244
rect 7232 21184 7296 21188
rect 10912 21244 10976 21248
rect 10912 21188 10916 21244
rect 10916 21188 10972 21244
rect 10972 21188 10976 21244
rect 10912 21184 10976 21188
rect 10992 21244 11056 21248
rect 10992 21188 10996 21244
rect 10996 21188 11052 21244
rect 11052 21188 11056 21244
rect 10992 21184 11056 21188
rect 11072 21244 11136 21248
rect 11072 21188 11076 21244
rect 11076 21188 11132 21244
rect 11132 21188 11136 21244
rect 11072 21184 11136 21188
rect 11152 21244 11216 21248
rect 11152 21188 11156 21244
rect 11156 21188 11212 21244
rect 11212 21188 11216 21244
rect 11152 21184 11216 21188
rect 11232 21244 11296 21248
rect 11232 21188 11236 21244
rect 11236 21188 11292 21244
rect 11292 21188 11296 21244
rect 11232 21184 11296 21188
rect 14912 21244 14976 21248
rect 14912 21188 14916 21244
rect 14916 21188 14972 21244
rect 14972 21188 14976 21244
rect 14912 21184 14976 21188
rect 14992 21244 15056 21248
rect 14992 21188 14996 21244
rect 14996 21188 15052 21244
rect 15052 21188 15056 21244
rect 14992 21184 15056 21188
rect 15072 21244 15136 21248
rect 15072 21188 15076 21244
rect 15076 21188 15132 21244
rect 15132 21188 15136 21244
rect 15072 21184 15136 21188
rect 15152 21244 15216 21248
rect 15152 21188 15156 21244
rect 15156 21188 15212 21244
rect 15212 21188 15216 21244
rect 15152 21184 15216 21188
rect 15232 21244 15296 21248
rect 15232 21188 15236 21244
rect 15236 21188 15292 21244
rect 15292 21188 15296 21244
rect 15232 21184 15296 21188
rect 18912 21244 18976 21248
rect 18912 21188 18916 21244
rect 18916 21188 18972 21244
rect 18972 21188 18976 21244
rect 18912 21184 18976 21188
rect 18992 21244 19056 21248
rect 18992 21188 18996 21244
rect 18996 21188 19052 21244
rect 19052 21188 19056 21244
rect 18992 21184 19056 21188
rect 19072 21244 19136 21248
rect 19072 21188 19076 21244
rect 19076 21188 19132 21244
rect 19132 21188 19136 21244
rect 19072 21184 19136 21188
rect 19152 21244 19216 21248
rect 19152 21188 19156 21244
rect 19156 21188 19212 21244
rect 19212 21188 19216 21244
rect 19152 21184 19216 21188
rect 19232 21244 19296 21248
rect 19232 21188 19236 21244
rect 19236 21188 19292 21244
rect 19292 21188 19296 21244
rect 19232 21184 19296 21188
rect 22912 21244 22976 21248
rect 22912 21188 22916 21244
rect 22916 21188 22972 21244
rect 22972 21188 22976 21244
rect 22912 21184 22976 21188
rect 22992 21244 23056 21248
rect 22992 21188 22996 21244
rect 22996 21188 23052 21244
rect 23052 21188 23056 21244
rect 22992 21184 23056 21188
rect 23072 21244 23136 21248
rect 23072 21188 23076 21244
rect 23076 21188 23132 21244
rect 23132 21188 23136 21244
rect 23072 21184 23136 21188
rect 23152 21244 23216 21248
rect 23152 21188 23156 21244
rect 23156 21188 23212 21244
rect 23212 21188 23216 21244
rect 23152 21184 23216 21188
rect 23232 21244 23296 21248
rect 23232 21188 23236 21244
rect 23236 21188 23292 21244
rect 23292 21188 23296 21244
rect 23232 21184 23296 21188
rect 19380 20844 19444 20908
rect 3652 20700 3716 20704
rect 3652 20644 3656 20700
rect 3656 20644 3712 20700
rect 3712 20644 3716 20700
rect 3652 20640 3716 20644
rect 3732 20700 3796 20704
rect 3732 20644 3736 20700
rect 3736 20644 3792 20700
rect 3792 20644 3796 20700
rect 3732 20640 3796 20644
rect 3812 20700 3876 20704
rect 3812 20644 3816 20700
rect 3816 20644 3872 20700
rect 3872 20644 3876 20700
rect 3812 20640 3876 20644
rect 3892 20700 3956 20704
rect 3892 20644 3896 20700
rect 3896 20644 3952 20700
rect 3952 20644 3956 20700
rect 3892 20640 3956 20644
rect 3972 20700 4036 20704
rect 3972 20644 3976 20700
rect 3976 20644 4032 20700
rect 4032 20644 4036 20700
rect 3972 20640 4036 20644
rect 7652 20700 7716 20704
rect 7652 20644 7656 20700
rect 7656 20644 7712 20700
rect 7712 20644 7716 20700
rect 7652 20640 7716 20644
rect 7732 20700 7796 20704
rect 7732 20644 7736 20700
rect 7736 20644 7792 20700
rect 7792 20644 7796 20700
rect 7732 20640 7796 20644
rect 7812 20700 7876 20704
rect 7812 20644 7816 20700
rect 7816 20644 7872 20700
rect 7872 20644 7876 20700
rect 7812 20640 7876 20644
rect 7892 20700 7956 20704
rect 7892 20644 7896 20700
rect 7896 20644 7952 20700
rect 7952 20644 7956 20700
rect 7892 20640 7956 20644
rect 7972 20700 8036 20704
rect 7972 20644 7976 20700
rect 7976 20644 8032 20700
rect 8032 20644 8036 20700
rect 7972 20640 8036 20644
rect 11652 20700 11716 20704
rect 11652 20644 11656 20700
rect 11656 20644 11712 20700
rect 11712 20644 11716 20700
rect 11652 20640 11716 20644
rect 11732 20700 11796 20704
rect 11732 20644 11736 20700
rect 11736 20644 11792 20700
rect 11792 20644 11796 20700
rect 11732 20640 11796 20644
rect 11812 20700 11876 20704
rect 11812 20644 11816 20700
rect 11816 20644 11872 20700
rect 11872 20644 11876 20700
rect 11812 20640 11876 20644
rect 11892 20700 11956 20704
rect 11892 20644 11896 20700
rect 11896 20644 11952 20700
rect 11952 20644 11956 20700
rect 11892 20640 11956 20644
rect 11972 20700 12036 20704
rect 11972 20644 11976 20700
rect 11976 20644 12032 20700
rect 12032 20644 12036 20700
rect 11972 20640 12036 20644
rect 15652 20700 15716 20704
rect 15652 20644 15656 20700
rect 15656 20644 15712 20700
rect 15712 20644 15716 20700
rect 15652 20640 15716 20644
rect 15732 20700 15796 20704
rect 15732 20644 15736 20700
rect 15736 20644 15792 20700
rect 15792 20644 15796 20700
rect 15732 20640 15796 20644
rect 15812 20700 15876 20704
rect 15812 20644 15816 20700
rect 15816 20644 15872 20700
rect 15872 20644 15876 20700
rect 15812 20640 15876 20644
rect 15892 20700 15956 20704
rect 15892 20644 15896 20700
rect 15896 20644 15952 20700
rect 15952 20644 15956 20700
rect 15892 20640 15956 20644
rect 15972 20700 16036 20704
rect 15972 20644 15976 20700
rect 15976 20644 16032 20700
rect 16032 20644 16036 20700
rect 15972 20640 16036 20644
rect 19652 20700 19716 20704
rect 19652 20644 19656 20700
rect 19656 20644 19712 20700
rect 19712 20644 19716 20700
rect 19652 20640 19716 20644
rect 19732 20700 19796 20704
rect 19732 20644 19736 20700
rect 19736 20644 19792 20700
rect 19792 20644 19796 20700
rect 19732 20640 19796 20644
rect 19812 20700 19876 20704
rect 19812 20644 19816 20700
rect 19816 20644 19872 20700
rect 19872 20644 19876 20700
rect 19812 20640 19876 20644
rect 19892 20700 19956 20704
rect 19892 20644 19896 20700
rect 19896 20644 19952 20700
rect 19952 20644 19956 20700
rect 19892 20640 19956 20644
rect 19972 20700 20036 20704
rect 19972 20644 19976 20700
rect 19976 20644 20032 20700
rect 20032 20644 20036 20700
rect 19972 20640 20036 20644
rect 23652 20700 23716 20704
rect 23652 20644 23656 20700
rect 23656 20644 23712 20700
rect 23712 20644 23716 20700
rect 23652 20640 23716 20644
rect 23732 20700 23796 20704
rect 23732 20644 23736 20700
rect 23736 20644 23792 20700
rect 23792 20644 23796 20700
rect 23732 20640 23796 20644
rect 23812 20700 23876 20704
rect 23812 20644 23816 20700
rect 23816 20644 23872 20700
rect 23872 20644 23876 20700
rect 23812 20640 23876 20644
rect 23892 20700 23956 20704
rect 23892 20644 23896 20700
rect 23896 20644 23952 20700
rect 23952 20644 23956 20700
rect 23892 20640 23956 20644
rect 23972 20700 24036 20704
rect 23972 20644 23976 20700
rect 23976 20644 24032 20700
rect 24032 20644 24036 20700
rect 23972 20640 24036 20644
rect 18276 20360 18340 20364
rect 18276 20304 18326 20360
rect 18326 20304 18340 20360
rect 18276 20300 18340 20304
rect 2912 20156 2976 20160
rect 2912 20100 2916 20156
rect 2916 20100 2972 20156
rect 2972 20100 2976 20156
rect 2912 20096 2976 20100
rect 2992 20156 3056 20160
rect 2992 20100 2996 20156
rect 2996 20100 3052 20156
rect 3052 20100 3056 20156
rect 2992 20096 3056 20100
rect 3072 20156 3136 20160
rect 3072 20100 3076 20156
rect 3076 20100 3132 20156
rect 3132 20100 3136 20156
rect 3072 20096 3136 20100
rect 3152 20156 3216 20160
rect 3152 20100 3156 20156
rect 3156 20100 3212 20156
rect 3212 20100 3216 20156
rect 3152 20096 3216 20100
rect 3232 20156 3296 20160
rect 3232 20100 3236 20156
rect 3236 20100 3292 20156
rect 3292 20100 3296 20156
rect 3232 20096 3296 20100
rect 6912 20156 6976 20160
rect 6912 20100 6916 20156
rect 6916 20100 6972 20156
rect 6972 20100 6976 20156
rect 6912 20096 6976 20100
rect 6992 20156 7056 20160
rect 6992 20100 6996 20156
rect 6996 20100 7052 20156
rect 7052 20100 7056 20156
rect 6992 20096 7056 20100
rect 7072 20156 7136 20160
rect 7072 20100 7076 20156
rect 7076 20100 7132 20156
rect 7132 20100 7136 20156
rect 7072 20096 7136 20100
rect 7152 20156 7216 20160
rect 7152 20100 7156 20156
rect 7156 20100 7212 20156
rect 7212 20100 7216 20156
rect 7152 20096 7216 20100
rect 7232 20156 7296 20160
rect 7232 20100 7236 20156
rect 7236 20100 7292 20156
rect 7292 20100 7296 20156
rect 7232 20096 7296 20100
rect 10912 20156 10976 20160
rect 10912 20100 10916 20156
rect 10916 20100 10972 20156
rect 10972 20100 10976 20156
rect 10912 20096 10976 20100
rect 10992 20156 11056 20160
rect 10992 20100 10996 20156
rect 10996 20100 11052 20156
rect 11052 20100 11056 20156
rect 10992 20096 11056 20100
rect 11072 20156 11136 20160
rect 11072 20100 11076 20156
rect 11076 20100 11132 20156
rect 11132 20100 11136 20156
rect 11072 20096 11136 20100
rect 11152 20156 11216 20160
rect 11152 20100 11156 20156
rect 11156 20100 11212 20156
rect 11212 20100 11216 20156
rect 11152 20096 11216 20100
rect 11232 20156 11296 20160
rect 11232 20100 11236 20156
rect 11236 20100 11292 20156
rect 11292 20100 11296 20156
rect 11232 20096 11296 20100
rect 14912 20156 14976 20160
rect 14912 20100 14916 20156
rect 14916 20100 14972 20156
rect 14972 20100 14976 20156
rect 14912 20096 14976 20100
rect 14992 20156 15056 20160
rect 14992 20100 14996 20156
rect 14996 20100 15052 20156
rect 15052 20100 15056 20156
rect 14992 20096 15056 20100
rect 15072 20156 15136 20160
rect 15072 20100 15076 20156
rect 15076 20100 15132 20156
rect 15132 20100 15136 20156
rect 15072 20096 15136 20100
rect 15152 20156 15216 20160
rect 15152 20100 15156 20156
rect 15156 20100 15212 20156
rect 15212 20100 15216 20156
rect 15152 20096 15216 20100
rect 15232 20156 15296 20160
rect 15232 20100 15236 20156
rect 15236 20100 15292 20156
rect 15292 20100 15296 20156
rect 15232 20096 15296 20100
rect 18912 20156 18976 20160
rect 18912 20100 18916 20156
rect 18916 20100 18972 20156
rect 18972 20100 18976 20156
rect 18912 20096 18976 20100
rect 18992 20156 19056 20160
rect 18992 20100 18996 20156
rect 18996 20100 19052 20156
rect 19052 20100 19056 20156
rect 18992 20096 19056 20100
rect 19072 20156 19136 20160
rect 19072 20100 19076 20156
rect 19076 20100 19132 20156
rect 19132 20100 19136 20156
rect 19072 20096 19136 20100
rect 19152 20156 19216 20160
rect 19152 20100 19156 20156
rect 19156 20100 19212 20156
rect 19212 20100 19216 20156
rect 19152 20096 19216 20100
rect 19232 20156 19296 20160
rect 19232 20100 19236 20156
rect 19236 20100 19292 20156
rect 19292 20100 19296 20156
rect 19232 20096 19296 20100
rect 22912 20156 22976 20160
rect 22912 20100 22916 20156
rect 22916 20100 22972 20156
rect 22972 20100 22976 20156
rect 22912 20096 22976 20100
rect 22992 20156 23056 20160
rect 22992 20100 22996 20156
rect 22996 20100 23052 20156
rect 23052 20100 23056 20156
rect 22992 20096 23056 20100
rect 23072 20156 23136 20160
rect 23072 20100 23076 20156
rect 23076 20100 23132 20156
rect 23132 20100 23136 20156
rect 23072 20096 23136 20100
rect 23152 20156 23216 20160
rect 23152 20100 23156 20156
rect 23156 20100 23212 20156
rect 23212 20100 23216 20156
rect 23152 20096 23216 20100
rect 23232 20156 23296 20160
rect 23232 20100 23236 20156
rect 23236 20100 23292 20156
rect 23292 20100 23296 20156
rect 23232 20096 23296 20100
rect 3652 19612 3716 19616
rect 3652 19556 3656 19612
rect 3656 19556 3712 19612
rect 3712 19556 3716 19612
rect 3652 19552 3716 19556
rect 3732 19612 3796 19616
rect 3732 19556 3736 19612
rect 3736 19556 3792 19612
rect 3792 19556 3796 19612
rect 3732 19552 3796 19556
rect 3812 19612 3876 19616
rect 3812 19556 3816 19612
rect 3816 19556 3872 19612
rect 3872 19556 3876 19612
rect 3812 19552 3876 19556
rect 3892 19612 3956 19616
rect 3892 19556 3896 19612
rect 3896 19556 3952 19612
rect 3952 19556 3956 19612
rect 3892 19552 3956 19556
rect 3972 19612 4036 19616
rect 3972 19556 3976 19612
rect 3976 19556 4032 19612
rect 4032 19556 4036 19612
rect 3972 19552 4036 19556
rect 7652 19612 7716 19616
rect 7652 19556 7656 19612
rect 7656 19556 7712 19612
rect 7712 19556 7716 19612
rect 7652 19552 7716 19556
rect 7732 19612 7796 19616
rect 7732 19556 7736 19612
rect 7736 19556 7792 19612
rect 7792 19556 7796 19612
rect 7732 19552 7796 19556
rect 7812 19612 7876 19616
rect 7812 19556 7816 19612
rect 7816 19556 7872 19612
rect 7872 19556 7876 19612
rect 7812 19552 7876 19556
rect 7892 19612 7956 19616
rect 7892 19556 7896 19612
rect 7896 19556 7952 19612
rect 7952 19556 7956 19612
rect 7892 19552 7956 19556
rect 7972 19612 8036 19616
rect 7972 19556 7976 19612
rect 7976 19556 8032 19612
rect 8032 19556 8036 19612
rect 7972 19552 8036 19556
rect 11652 19612 11716 19616
rect 11652 19556 11656 19612
rect 11656 19556 11712 19612
rect 11712 19556 11716 19612
rect 11652 19552 11716 19556
rect 11732 19612 11796 19616
rect 11732 19556 11736 19612
rect 11736 19556 11792 19612
rect 11792 19556 11796 19612
rect 11732 19552 11796 19556
rect 11812 19612 11876 19616
rect 11812 19556 11816 19612
rect 11816 19556 11872 19612
rect 11872 19556 11876 19612
rect 11812 19552 11876 19556
rect 11892 19612 11956 19616
rect 11892 19556 11896 19612
rect 11896 19556 11952 19612
rect 11952 19556 11956 19612
rect 11892 19552 11956 19556
rect 11972 19612 12036 19616
rect 11972 19556 11976 19612
rect 11976 19556 12032 19612
rect 12032 19556 12036 19612
rect 11972 19552 12036 19556
rect 15652 19612 15716 19616
rect 15652 19556 15656 19612
rect 15656 19556 15712 19612
rect 15712 19556 15716 19612
rect 15652 19552 15716 19556
rect 15732 19612 15796 19616
rect 15732 19556 15736 19612
rect 15736 19556 15792 19612
rect 15792 19556 15796 19612
rect 15732 19552 15796 19556
rect 15812 19612 15876 19616
rect 15812 19556 15816 19612
rect 15816 19556 15872 19612
rect 15872 19556 15876 19612
rect 15812 19552 15876 19556
rect 15892 19612 15956 19616
rect 15892 19556 15896 19612
rect 15896 19556 15952 19612
rect 15952 19556 15956 19612
rect 15892 19552 15956 19556
rect 15972 19612 16036 19616
rect 15972 19556 15976 19612
rect 15976 19556 16032 19612
rect 16032 19556 16036 19612
rect 15972 19552 16036 19556
rect 19652 19612 19716 19616
rect 19652 19556 19656 19612
rect 19656 19556 19712 19612
rect 19712 19556 19716 19612
rect 19652 19552 19716 19556
rect 19732 19612 19796 19616
rect 19732 19556 19736 19612
rect 19736 19556 19792 19612
rect 19792 19556 19796 19612
rect 19732 19552 19796 19556
rect 19812 19612 19876 19616
rect 19812 19556 19816 19612
rect 19816 19556 19872 19612
rect 19872 19556 19876 19612
rect 19812 19552 19876 19556
rect 19892 19612 19956 19616
rect 19892 19556 19896 19612
rect 19896 19556 19952 19612
rect 19952 19556 19956 19612
rect 19892 19552 19956 19556
rect 19972 19612 20036 19616
rect 19972 19556 19976 19612
rect 19976 19556 20032 19612
rect 20032 19556 20036 19612
rect 19972 19552 20036 19556
rect 23652 19612 23716 19616
rect 23652 19556 23656 19612
rect 23656 19556 23712 19612
rect 23712 19556 23716 19612
rect 23652 19552 23716 19556
rect 23732 19612 23796 19616
rect 23732 19556 23736 19612
rect 23736 19556 23792 19612
rect 23792 19556 23796 19612
rect 23732 19552 23796 19556
rect 23812 19612 23876 19616
rect 23812 19556 23816 19612
rect 23816 19556 23872 19612
rect 23872 19556 23876 19612
rect 23812 19552 23876 19556
rect 23892 19612 23956 19616
rect 23892 19556 23896 19612
rect 23896 19556 23952 19612
rect 23952 19556 23956 19612
rect 23892 19552 23956 19556
rect 23972 19612 24036 19616
rect 23972 19556 23976 19612
rect 23976 19556 24032 19612
rect 24032 19556 24036 19612
rect 23972 19552 24036 19556
rect 5212 19408 5276 19412
rect 5212 19352 5262 19408
rect 5262 19352 5276 19408
rect 5212 19348 5276 19352
rect 9996 19212 10060 19276
rect 2912 19068 2976 19072
rect 2912 19012 2916 19068
rect 2916 19012 2972 19068
rect 2972 19012 2976 19068
rect 2912 19008 2976 19012
rect 2992 19068 3056 19072
rect 2992 19012 2996 19068
rect 2996 19012 3052 19068
rect 3052 19012 3056 19068
rect 2992 19008 3056 19012
rect 3072 19068 3136 19072
rect 3072 19012 3076 19068
rect 3076 19012 3132 19068
rect 3132 19012 3136 19068
rect 3072 19008 3136 19012
rect 3152 19068 3216 19072
rect 3152 19012 3156 19068
rect 3156 19012 3212 19068
rect 3212 19012 3216 19068
rect 3152 19008 3216 19012
rect 3232 19068 3296 19072
rect 3232 19012 3236 19068
rect 3236 19012 3292 19068
rect 3292 19012 3296 19068
rect 3232 19008 3296 19012
rect 6912 19068 6976 19072
rect 6912 19012 6916 19068
rect 6916 19012 6972 19068
rect 6972 19012 6976 19068
rect 6912 19008 6976 19012
rect 6992 19068 7056 19072
rect 6992 19012 6996 19068
rect 6996 19012 7052 19068
rect 7052 19012 7056 19068
rect 6992 19008 7056 19012
rect 7072 19068 7136 19072
rect 7072 19012 7076 19068
rect 7076 19012 7132 19068
rect 7132 19012 7136 19068
rect 7072 19008 7136 19012
rect 7152 19068 7216 19072
rect 7152 19012 7156 19068
rect 7156 19012 7212 19068
rect 7212 19012 7216 19068
rect 7152 19008 7216 19012
rect 7232 19068 7296 19072
rect 7232 19012 7236 19068
rect 7236 19012 7292 19068
rect 7292 19012 7296 19068
rect 7232 19008 7296 19012
rect 10912 19068 10976 19072
rect 10912 19012 10916 19068
rect 10916 19012 10972 19068
rect 10972 19012 10976 19068
rect 10912 19008 10976 19012
rect 10992 19068 11056 19072
rect 10992 19012 10996 19068
rect 10996 19012 11052 19068
rect 11052 19012 11056 19068
rect 10992 19008 11056 19012
rect 11072 19068 11136 19072
rect 11072 19012 11076 19068
rect 11076 19012 11132 19068
rect 11132 19012 11136 19068
rect 11072 19008 11136 19012
rect 11152 19068 11216 19072
rect 11152 19012 11156 19068
rect 11156 19012 11212 19068
rect 11212 19012 11216 19068
rect 11152 19008 11216 19012
rect 11232 19068 11296 19072
rect 11232 19012 11236 19068
rect 11236 19012 11292 19068
rect 11292 19012 11296 19068
rect 11232 19008 11296 19012
rect 14912 19068 14976 19072
rect 14912 19012 14916 19068
rect 14916 19012 14972 19068
rect 14972 19012 14976 19068
rect 14912 19008 14976 19012
rect 14992 19068 15056 19072
rect 14992 19012 14996 19068
rect 14996 19012 15052 19068
rect 15052 19012 15056 19068
rect 14992 19008 15056 19012
rect 15072 19068 15136 19072
rect 15072 19012 15076 19068
rect 15076 19012 15132 19068
rect 15132 19012 15136 19068
rect 15072 19008 15136 19012
rect 15152 19068 15216 19072
rect 15152 19012 15156 19068
rect 15156 19012 15212 19068
rect 15212 19012 15216 19068
rect 15152 19008 15216 19012
rect 15232 19068 15296 19072
rect 15232 19012 15236 19068
rect 15236 19012 15292 19068
rect 15292 19012 15296 19068
rect 15232 19008 15296 19012
rect 18912 19068 18976 19072
rect 18912 19012 18916 19068
rect 18916 19012 18972 19068
rect 18972 19012 18976 19068
rect 18912 19008 18976 19012
rect 18992 19068 19056 19072
rect 18992 19012 18996 19068
rect 18996 19012 19052 19068
rect 19052 19012 19056 19068
rect 18992 19008 19056 19012
rect 19072 19068 19136 19072
rect 19072 19012 19076 19068
rect 19076 19012 19132 19068
rect 19132 19012 19136 19068
rect 19072 19008 19136 19012
rect 19152 19068 19216 19072
rect 19152 19012 19156 19068
rect 19156 19012 19212 19068
rect 19212 19012 19216 19068
rect 19152 19008 19216 19012
rect 19232 19068 19296 19072
rect 19232 19012 19236 19068
rect 19236 19012 19292 19068
rect 19292 19012 19296 19068
rect 19232 19008 19296 19012
rect 22912 19068 22976 19072
rect 22912 19012 22916 19068
rect 22916 19012 22972 19068
rect 22972 19012 22976 19068
rect 22912 19008 22976 19012
rect 22992 19068 23056 19072
rect 22992 19012 22996 19068
rect 22996 19012 23052 19068
rect 23052 19012 23056 19068
rect 22992 19008 23056 19012
rect 23072 19068 23136 19072
rect 23072 19012 23076 19068
rect 23076 19012 23132 19068
rect 23132 19012 23136 19068
rect 23072 19008 23136 19012
rect 23152 19068 23216 19072
rect 23152 19012 23156 19068
rect 23156 19012 23212 19068
rect 23212 19012 23216 19068
rect 23152 19008 23216 19012
rect 23232 19068 23296 19072
rect 23232 19012 23236 19068
rect 23236 19012 23292 19068
rect 23292 19012 23296 19068
rect 23232 19008 23296 19012
rect 3652 18524 3716 18528
rect 3652 18468 3656 18524
rect 3656 18468 3712 18524
rect 3712 18468 3716 18524
rect 3652 18464 3716 18468
rect 3732 18524 3796 18528
rect 3732 18468 3736 18524
rect 3736 18468 3792 18524
rect 3792 18468 3796 18524
rect 3732 18464 3796 18468
rect 3812 18524 3876 18528
rect 3812 18468 3816 18524
rect 3816 18468 3872 18524
rect 3872 18468 3876 18524
rect 3812 18464 3876 18468
rect 3892 18524 3956 18528
rect 3892 18468 3896 18524
rect 3896 18468 3952 18524
rect 3952 18468 3956 18524
rect 3892 18464 3956 18468
rect 3972 18524 4036 18528
rect 3972 18468 3976 18524
rect 3976 18468 4032 18524
rect 4032 18468 4036 18524
rect 3972 18464 4036 18468
rect 7652 18524 7716 18528
rect 7652 18468 7656 18524
rect 7656 18468 7712 18524
rect 7712 18468 7716 18524
rect 7652 18464 7716 18468
rect 7732 18524 7796 18528
rect 7732 18468 7736 18524
rect 7736 18468 7792 18524
rect 7792 18468 7796 18524
rect 7732 18464 7796 18468
rect 7812 18524 7876 18528
rect 7812 18468 7816 18524
rect 7816 18468 7872 18524
rect 7872 18468 7876 18524
rect 7812 18464 7876 18468
rect 7892 18524 7956 18528
rect 7892 18468 7896 18524
rect 7896 18468 7952 18524
rect 7952 18468 7956 18524
rect 7892 18464 7956 18468
rect 7972 18524 8036 18528
rect 7972 18468 7976 18524
rect 7976 18468 8032 18524
rect 8032 18468 8036 18524
rect 7972 18464 8036 18468
rect 11652 18524 11716 18528
rect 11652 18468 11656 18524
rect 11656 18468 11712 18524
rect 11712 18468 11716 18524
rect 11652 18464 11716 18468
rect 11732 18524 11796 18528
rect 11732 18468 11736 18524
rect 11736 18468 11792 18524
rect 11792 18468 11796 18524
rect 11732 18464 11796 18468
rect 11812 18524 11876 18528
rect 11812 18468 11816 18524
rect 11816 18468 11872 18524
rect 11872 18468 11876 18524
rect 11812 18464 11876 18468
rect 11892 18524 11956 18528
rect 11892 18468 11896 18524
rect 11896 18468 11952 18524
rect 11952 18468 11956 18524
rect 11892 18464 11956 18468
rect 11972 18524 12036 18528
rect 11972 18468 11976 18524
rect 11976 18468 12032 18524
rect 12032 18468 12036 18524
rect 11972 18464 12036 18468
rect 15652 18524 15716 18528
rect 15652 18468 15656 18524
rect 15656 18468 15712 18524
rect 15712 18468 15716 18524
rect 15652 18464 15716 18468
rect 15732 18524 15796 18528
rect 15732 18468 15736 18524
rect 15736 18468 15792 18524
rect 15792 18468 15796 18524
rect 15732 18464 15796 18468
rect 15812 18524 15876 18528
rect 15812 18468 15816 18524
rect 15816 18468 15872 18524
rect 15872 18468 15876 18524
rect 15812 18464 15876 18468
rect 15892 18524 15956 18528
rect 15892 18468 15896 18524
rect 15896 18468 15952 18524
rect 15952 18468 15956 18524
rect 15892 18464 15956 18468
rect 15972 18524 16036 18528
rect 15972 18468 15976 18524
rect 15976 18468 16032 18524
rect 16032 18468 16036 18524
rect 15972 18464 16036 18468
rect 19652 18524 19716 18528
rect 19652 18468 19656 18524
rect 19656 18468 19712 18524
rect 19712 18468 19716 18524
rect 19652 18464 19716 18468
rect 19732 18524 19796 18528
rect 19732 18468 19736 18524
rect 19736 18468 19792 18524
rect 19792 18468 19796 18524
rect 19732 18464 19796 18468
rect 19812 18524 19876 18528
rect 19812 18468 19816 18524
rect 19816 18468 19872 18524
rect 19872 18468 19876 18524
rect 19812 18464 19876 18468
rect 19892 18524 19956 18528
rect 19892 18468 19896 18524
rect 19896 18468 19952 18524
rect 19952 18468 19956 18524
rect 19892 18464 19956 18468
rect 19972 18524 20036 18528
rect 19972 18468 19976 18524
rect 19976 18468 20032 18524
rect 20032 18468 20036 18524
rect 19972 18464 20036 18468
rect 23652 18524 23716 18528
rect 23652 18468 23656 18524
rect 23656 18468 23712 18524
rect 23712 18468 23716 18524
rect 23652 18464 23716 18468
rect 23732 18524 23796 18528
rect 23732 18468 23736 18524
rect 23736 18468 23792 18524
rect 23792 18468 23796 18524
rect 23732 18464 23796 18468
rect 23812 18524 23876 18528
rect 23812 18468 23816 18524
rect 23816 18468 23872 18524
rect 23872 18468 23876 18524
rect 23812 18464 23876 18468
rect 23892 18524 23956 18528
rect 23892 18468 23896 18524
rect 23896 18468 23952 18524
rect 23952 18468 23956 18524
rect 23892 18464 23956 18468
rect 23972 18524 24036 18528
rect 23972 18468 23976 18524
rect 23976 18468 24032 18524
rect 24032 18468 24036 18524
rect 23972 18464 24036 18468
rect 14596 18124 14660 18188
rect 2912 17980 2976 17984
rect 2912 17924 2916 17980
rect 2916 17924 2972 17980
rect 2972 17924 2976 17980
rect 2912 17920 2976 17924
rect 2992 17980 3056 17984
rect 2992 17924 2996 17980
rect 2996 17924 3052 17980
rect 3052 17924 3056 17980
rect 2992 17920 3056 17924
rect 3072 17980 3136 17984
rect 3072 17924 3076 17980
rect 3076 17924 3132 17980
rect 3132 17924 3136 17980
rect 3072 17920 3136 17924
rect 3152 17980 3216 17984
rect 3152 17924 3156 17980
rect 3156 17924 3212 17980
rect 3212 17924 3216 17980
rect 3152 17920 3216 17924
rect 3232 17980 3296 17984
rect 3232 17924 3236 17980
rect 3236 17924 3292 17980
rect 3292 17924 3296 17980
rect 3232 17920 3296 17924
rect 6912 17980 6976 17984
rect 6912 17924 6916 17980
rect 6916 17924 6972 17980
rect 6972 17924 6976 17980
rect 6912 17920 6976 17924
rect 6992 17980 7056 17984
rect 6992 17924 6996 17980
rect 6996 17924 7052 17980
rect 7052 17924 7056 17980
rect 6992 17920 7056 17924
rect 7072 17980 7136 17984
rect 7072 17924 7076 17980
rect 7076 17924 7132 17980
rect 7132 17924 7136 17980
rect 7072 17920 7136 17924
rect 7152 17980 7216 17984
rect 7152 17924 7156 17980
rect 7156 17924 7212 17980
rect 7212 17924 7216 17980
rect 7152 17920 7216 17924
rect 7232 17980 7296 17984
rect 7232 17924 7236 17980
rect 7236 17924 7292 17980
rect 7292 17924 7296 17980
rect 7232 17920 7296 17924
rect 10912 17980 10976 17984
rect 10912 17924 10916 17980
rect 10916 17924 10972 17980
rect 10972 17924 10976 17980
rect 10912 17920 10976 17924
rect 10992 17980 11056 17984
rect 10992 17924 10996 17980
rect 10996 17924 11052 17980
rect 11052 17924 11056 17980
rect 10992 17920 11056 17924
rect 11072 17980 11136 17984
rect 11072 17924 11076 17980
rect 11076 17924 11132 17980
rect 11132 17924 11136 17980
rect 11072 17920 11136 17924
rect 11152 17980 11216 17984
rect 11152 17924 11156 17980
rect 11156 17924 11212 17980
rect 11212 17924 11216 17980
rect 11152 17920 11216 17924
rect 11232 17980 11296 17984
rect 11232 17924 11236 17980
rect 11236 17924 11292 17980
rect 11292 17924 11296 17980
rect 11232 17920 11296 17924
rect 14912 17980 14976 17984
rect 14912 17924 14916 17980
rect 14916 17924 14972 17980
rect 14972 17924 14976 17980
rect 14912 17920 14976 17924
rect 14992 17980 15056 17984
rect 14992 17924 14996 17980
rect 14996 17924 15052 17980
rect 15052 17924 15056 17980
rect 14992 17920 15056 17924
rect 15072 17980 15136 17984
rect 15072 17924 15076 17980
rect 15076 17924 15132 17980
rect 15132 17924 15136 17980
rect 15072 17920 15136 17924
rect 15152 17980 15216 17984
rect 15152 17924 15156 17980
rect 15156 17924 15212 17980
rect 15212 17924 15216 17980
rect 15152 17920 15216 17924
rect 15232 17980 15296 17984
rect 15232 17924 15236 17980
rect 15236 17924 15292 17980
rect 15292 17924 15296 17980
rect 15232 17920 15296 17924
rect 18912 17980 18976 17984
rect 18912 17924 18916 17980
rect 18916 17924 18972 17980
rect 18972 17924 18976 17980
rect 18912 17920 18976 17924
rect 18992 17980 19056 17984
rect 18992 17924 18996 17980
rect 18996 17924 19052 17980
rect 19052 17924 19056 17980
rect 18992 17920 19056 17924
rect 19072 17980 19136 17984
rect 19072 17924 19076 17980
rect 19076 17924 19132 17980
rect 19132 17924 19136 17980
rect 19072 17920 19136 17924
rect 19152 17980 19216 17984
rect 19152 17924 19156 17980
rect 19156 17924 19212 17980
rect 19212 17924 19216 17980
rect 19152 17920 19216 17924
rect 19232 17980 19296 17984
rect 19232 17924 19236 17980
rect 19236 17924 19292 17980
rect 19292 17924 19296 17980
rect 19232 17920 19296 17924
rect 22912 17980 22976 17984
rect 22912 17924 22916 17980
rect 22916 17924 22972 17980
rect 22972 17924 22976 17980
rect 22912 17920 22976 17924
rect 22992 17980 23056 17984
rect 22992 17924 22996 17980
rect 22996 17924 23052 17980
rect 23052 17924 23056 17980
rect 22992 17920 23056 17924
rect 23072 17980 23136 17984
rect 23072 17924 23076 17980
rect 23076 17924 23132 17980
rect 23132 17924 23136 17980
rect 23072 17920 23136 17924
rect 23152 17980 23216 17984
rect 23152 17924 23156 17980
rect 23156 17924 23212 17980
rect 23212 17924 23216 17980
rect 23152 17920 23216 17924
rect 23232 17980 23296 17984
rect 23232 17924 23236 17980
rect 23236 17924 23292 17980
rect 23292 17924 23296 17980
rect 23232 17920 23296 17924
rect 3652 17436 3716 17440
rect 3652 17380 3656 17436
rect 3656 17380 3712 17436
rect 3712 17380 3716 17436
rect 3652 17376 3716 17380
rect 3732 17436 3796 17440
rect 3732 17380 3736 17436
rect 3736 17380 3792 17436
rect 3792 17380 3796 17436
rect 3732 17376 3796 17380
rect 3812 17436 3876 17440
rect 3812 17380 3816 17436
rect 3816 17380 3872 17436
rect 3872 17380 3876 17436
rect 3812 17376 3876 17380
rect 3892 17436 3956 17440
rect 3892 17380 3896 17436
rect 3896 17380 3952 17436
rect 3952 17380 3956 17436
rect 3892 17376 3956 17380
rect 3972 17436 4036 17440
rect 3972 17380 3976 17436
rect 3976 17380 4032 17436
rect 4032 17380 4036 17436
rect 3972 17376 4036 17380
rect 7652 17436 7716 17440
rect 7652 17380 7656 17436
rect 7656 17380 7712 17436
rect 7712 17380 7716 17436
rect 7652 17376 7716 17380
rect 7732 17436 7796 17440
rect 7732 17380 7736 17436
rect 7736 17380 7792 17436
rect 7792 17380 7796 17436
rect 7732 17376 7796 17380
rect 7812 17436 7876 17440
rect 7812 17380 7816 17436
rect 7816 17380 7872 17436
rect 7872 17380 7876 17436
rect 7812 17376 7876 17380
rect 7892 17436 7956 17440
rect 7892 17380 7896 17436
rect 7896 17380 7952 17436
rect 7952 17380 7956 17436
rect 7892 17376 7956 17380
rect 7972 17436 8036 17440
rect 7972 17380 7976 17436
rect 7976 17380 8032 17436
rect 8032 17380 8036 17436
rect 7972 17376 8036 17380
rect 11652 17436 11716 17440
rect 11652 17380 11656 17436
rect 11656 17380 11712 17436
rect 11712 17380 11716 17436
rect 11652 17376 11716 17380
rect 11732 17436 11796 17440
rect 11732 17380 11736 17436
rect 11736 17380 11792 17436
rect 11792 17380 11796 17436
rect 11732 17376 11796 17380
rect 11812 17436 11876 17440
rect 11812 17380 11816 17436
rect 11816 17380 11872 17436
rect 11872 17380 11876 17436
rect 11812 17376 11876 17380
rect 11892 17436 11956 17440
rect 11892 17380 11896 17436
rect 11896 17380 11952 17436
rect 11952 17380 11956 17436
rect 11892 17376 11956 17380
rect 11972 17436 12036 17440
rect 11972 17380 11976 17436
rect 11976 17380 12032 17436
rect 12032 17380 12036 17436
rect 11972 17376 12036 17380
rect 15652 17436 15716 17440
rect 15652 17380 15656 17436
rect 15656 17380 15712 17436
rect 15712 17380 15716 17436
rect 15652 17376 15716 17380
rect 15732 17436 15796 17440
rect 15732 17380 15736 17436
rect 15736 17380 15792 17436
rect 15792 17380 15796 17436
rect 15732 17376 15796 17380
rect 15812 17436 15876 17440
rect 15812 17380 15816 17436
rect 15816 17380 15872 17436
rect 15872 17380 15876 17436
rect 15812 17376 15876 17380
rect 15892 17436 15956 17440
rect 15892 17380 15896 17436
rect 15896 17380 15952 17436
rect 15952 17380 15956 17436
rect 15892 17376 15956 17380
rect 15972 17436 16036 17440
rect 15972 17380 15976 17436
rect 15976 17380 16032 17436
rect 16032 17380 16036 17436
rect 15972 17376 16036 17380
rect 19652 17436 19716 17440
rect 19652 17380 19656 17436
rect 19656 17380 19712 17436
rect 19712 17380 19716 17436
rect 19652 17376 19716 17380
rect 19732 17436 19796 17440
rect 19732 17380 19736 17436
rect 19736 17380 19792 17436
rect 19792 17380 19796 17436
rect 19732 17376 19796 17380
rect 19812 17436 19876 17440
rect 19812 17380 19816 17436
rect 19816 17380 19872 17436
rect 19872 17380 19876 17436
rect 19812 17376 19876 17380
rect 19892 17436 19956 17440
rect 19892 17380 19896 17436
rect 19896 17380 19952 17436
rect 19952 17380 19956 17436
rect 19892 17376 19956 17380
rect 19972 17436 20036 17440
rect 19972 17380 19976 17436
rect 19976 17380 20032 17436
rect 20032 17380 20036 17436
rect 19972 17376 20036 17380
rect 23652 17436 23716 17440
rect 23652 17380 23656 17436
rect 23656 17380 23712 17436
rect 23712 17380 23716 17436
rect 23652 17376 23716 17380
rect 23732 17436 23796 17440
rect 23732 17380 23736 17436
rect 23736 17380 23792 17436
rect 23792 17380 23796 17436
rect 23732 17376 23796 17380
rect 23812 17436 23876 17440
rect 23812 17380 23816 17436
rect 23816 17380 23872 17436
rect 23872 17380 23876 17436
rect 23812 17376 23876 17380
rect 23892 17436 23956 17440
rect 23892 17380 23896 17436
rect 23896 17380 23952 17436
rect 23952 17380 23956 17436
rect 23892 17376 23956 17380
rect 23972 17436 24036 17440
rect 23972 17380 23976 17436
rect 23976 17380 24032 17436
rect 24032 17380 24036 17436
rect 23972 17376 24036 17380
rect 2912 16892 2976 16896
rect 2912 16836 2916 16892
rect 2916 16836 2972 16892
rect 2972 16836 2976 16892
rect 2912 16832 2976 16836
rect 2992 16892 3056 16896
rect 2992 16836 2996 16892
rect 2996 16836 3052 16892
rect 3052 16836 3056 16892
rect 2992 16832 3056 16836
rect 3072 16892 3136 16896
rect 3072 16836 3076 16892
rect 3076 16836 3132 16892
rect 3132 16836 3136 16892
rect 3072 16832 3136 16836
rect 3152 16892 3216 16896
rect 3152 16836 3156 16892
rect 3156 16836 3212 16892
rect 3212 16836 3216 16892
rect 3152 16832 3216 16836
rect 3232 16892 3296 16896
rect 3232 16836 3236 16892
rect 3236 16836 3292 16892
rect 3292 16836 3296 16892
rect 3232 16832 3296 16836
rect 6912 16892 6976 16896
rect 6912 16836 6916 16892
rect 6916 16836 6972 16892
rect 6972 16836 6976 16892
rect 6912 16832 6976 16836
rect 6992 16892 7056 16896
rect 6992 16836 6996 16892
rect 6996 16836 7052 16892
rect 7052 16836 7056 16892
rect 6992 16832 7056 16836
rect 7072 16892 7136 16896
rect 7072 16836 7076 16892
rect 7076 16836 7132 16892
rect 7132 16836 7136 16892
rect 7072 16832 7136 16836
rect 7152 16892 7216 16896
rect 7152 16836 7156 16892
rect 7156 16836 7212 16892
rect 7212 16836 7216 16892
rect 7152 16832 7216 16836
rect 7232 16892 7296 16896
rect 7232 16836 7236 16892
rect 7236 16836 7292 16892
rect 7292 16836 7296 16892
rect 7232 16832 7296 16836
rect 10912 16892 10976 16896
rect 10912 16836 10916 16892
rect 10916 16836 10972 16892
rect 10972 16836 10976 16892
rect 10912 16832 10976 16836
rect 10992 16892 11056 16896
rect 10992 16836 10996 16892
rect 10996 16836 11052 16892
rect 11052 16836 11056 16892
rect 10992 16832 11056 16836
rect 11072 16892 11136 16896
rect 11072 16836 11076 16892
rect 11076 16836 11132 16892
rect 11132 16836 11136 16892
rect 11072 16832 11136 16836
rect 11152 16892 11216 16896
rect 11152 16836 11156 16892
rect 11156 16836 11212 16892
rect 11212 16836 11216 16892
rect 11152 16832 11216 16836
rect 11232 16892 11296 16896
rect 11232 16836 11236 16892
rect 11236 16836 11292 16892
rect 11292 16836 11296 16892
rect 11232 16832 11296 16836
rect 14912 16892 14976 16896
rect 14912 16836 14916 16892
rect 14916 16836 14972 16892
rect 14972 16836 14976 16892
rect 14912 16832 14976 16836
rect 14992 16892 15056 16896
rect 14992 16836 14996 16892
rect 14996 16836 15052 16892
rect 15052 16836 15056 16892
rect 14992 16832 15056 16836
rect 15072 16892 15136 16896
rect 15072 16836 15076 16892
rect 15076 16836 15132 16892
rect 15132 16836 15136 16892
rect 15072 16832 15136 16836
rect 15152 16892 15216 16896
rect 15152 16836 15156 16892
rect 15156 16836 15212 16892
rect 15212 16836 15216 16892
rect 15152 16832 15216 16836
rect 15232 16892 15296 16896
rect 15232 16836 15236 16892
rect 15236 16836 15292 16892
rect 15292 16836 15296 16892
rect 15232 16832 15296 16836
rect 18912 16892 18976 16896
rect 18912 16836 18916 16892
rect 18916 16836 18972 16892
rect 18972 16836 18976 16892
rect 18912 16832 18976 16836
rect 18992 16892 19056 16896
rect 18992 16836 18996 16892
rect 18996 16836 19052 16892
rect 19052 16836 19056 16892
rect 18992 16832 19056 16836
rect 19072 16892 19136 16896
rect 19072 16836 19076 16892
rect 19076 16836 19132 16892
rect 19132 16836 19136 16892
rect 19072 16832 19136 16836
rect 19152 16892 19216 16896
rect 19152 16836 19156 16892
rect 19156 16836 19212 16892
rect 19212 16836 19216 16892
rect 19152 16832 19216 16836
rect 19232 16892 19296 16896
rect 19232 16836 19236 16892
rect 19236 16836 19292 16892
rect 19292 16836 19296 16892
rect 19232 16832 19296 16836
rect 22912 16892 22976 16896
rect 22912 16836 22916 16892
rect 22916 16836 22972 16892
rect 22972 16836 22976 16892
rect 22912 16832 22976 16836
rect 22992 16892 23056 16896
rect 22992 16836 22996 16892
rect 22996 16836 23052 16892
rect 23052 16836 23056 16892
rect 22992 16832 23056 16836
rect 23072 16892 23136 16896
rect 23072 16836 23076 16892
rect 23076 16836 23132 16892
rect 23132 16836 23136 16892
rect 23072 16832 23136 16836
rect 23152 16892 23216 16896
rect 23152 16836 23156 16892
rect 23156 16836 23212 16892
rect 23212 16836 23216 16892
rect 23152 16832 23216 16836
rect 23232 16892 23296 16896
rect 23232 16836 23236 16892
rect 23236 16836 23292 16892
rect 23292 16836 23296 16892
rect 23232 16832 23296 16836
rect 15516 16688 15580 16692
rect 15516 16632 15566 16688
rect 15566 16632 15580 16688
rect 15516 16628 15580 16632
rect 3652 16348 3716 16352
rect 3652 16292 3656 16348
rect 3656 16292 3712 16348
rect 3712 16292 3716 16348
rect 3652 16288 3716 16292
rect 3732 16348 3796 16352
rect 3732 16292 3736 16348
rect 3736 16292 3792 16348
rect 3792 16292 3796 16348
rect 3732 16288 3796 16292
rect 3812 16348 3876 16352
rect 3812 16292 3816 16348
rect 3816 16292 3872 16348
rect 3872 16292 3876 16348
rect 3812 16288 3876 16292
rect 3892 16348 3956 16352
rect 3892 16292 3896 16348
rect 3896 16292 3952 16348
rect 3952 16292 3956 16348
rect 3892 16288 3956 16292
rect 3972 16348 4036 16352
rect 3972 16292 3976 16348
rect 3976 16292 4032 16348
rect 4032 16292 4036 16348
rect 3972 16288 4036 16292
rect 7652 16348 7716 16352
rect 7652 16292 7656 16348
rect 7656 16292 7712 16348
rect 7712 16292 7716 16348
rect 7652 16288 7716 16292
rect 7732 16348 7796 16352
rect 7732 16292 7736 16348
rect 7736 16292 7792 16348
rect 7792 16292 7796 16348
rect 7732 16288 7796 16292
rect 7812 16348 7876 16352
rect 7812 16292 7816 16348
rect 7816 16292 7872 16348
rect 7872 16292 7876 16348
rect 7812 16288 7876 16292
rect 7892 16348 7956 16352
rect 7892 16292 7896 16348
rect 7896 16292 7952 16348
rect 7952 16292 7956 16348
rect 7892 16288 7956 16292
rect 7972 16348 8036 16352
rect 7972 16292 7976 16348
rect 7976 16292 8032 16348
rect 8032 16292 8036 16348
rect 7972 16288 8036 16292
rect 11652 16348 11716 16352
rect 11652 16292 11656 16348
rect 11656 16292 11712 16348
rect 11712 16292 11716 16348
rect 11652 16288 11716 16292
rect 11732 16348 11796 16352
rect 11732 16292 11736 16348
rect 11736 16292 11792 16348
rect 11792 16292 11796 16348
rect 11732 16288 11796 16292
rect 11812 16348 11876 16352
rect 11812 16292 11816 16348
rect 11816 16292 11872 16348
rect 11872 16292 11876 16348
rect 11812 16288 11876 16292
rect 11892 16348 11956 16352
rect 11892 16292 11896 16348
rect 11896 16292 11952 16348
rect 11952 16292 11956 16348
rect 11892 16288 11956 16292
rect 11972 16348 12036 16352
rect 11972 16292 11976 16348
rect 11976 16292 12032 16348
rect 12032 16292 12036 16348
rect 11972 16288 12036 16292
rect 15652 16348 15716 16352
rect 15652 16292 15656 16348
rect 15656 16292 15712 16348
rect 15712 16292 15716 16348
rect 15652 16288 15716 16292
rect 15732 16348 15796 16352
rect 15732 16292 15736 16348
rect 15736 16292 15792 16348
rect 15792 16292 15796 16348
rect 15732 16288 15796 16292
rect 15812 16348 15876 16352
rect 15812 16292 15816 16348
rect 15816 16292 15872 16348
rect 15872 16292 15876 16348
rect 15812 16288 15876 16292
rect 15892 16348 15956 16352
rect 15892 16292 15896 16348
rect 15896 16292 15952 16348
rect 15952 16292 15956 16348
rect 15892 16288 15956 16292
rect 15972 16348 16036 16352
rect 15972 16292 15976 16348
rect 15976 16292 16032 16348
rect 16032 16292 16036 16348
rect 15972 16288 16036 16292
rect 19652 16348 19716 16352
rect 19652 16292 19656 16348
rect 19656 16292 19712 16348
rect 19712 16292 19716 16348
rect 19652 16288 19716 16292
rect 19732 16348 19796 16352
rect 19732 16292 19736 16348
rect 19736 16292 19792 16348
rect 19792 16292 19796 16348
rect 19732 16288 19796 16292
rect 19812 16348 19876 16352
rect 19812 16292 19816 16348
rect 19816 16292 19872 16348
rect 19872 16292 19876 16348
rect 19812 16288 19876 16292
rect 19892 16348 19956 16352
rect 19892 16292 19896 16348
rect 19896 16292 19952 16348
rect 19952 16292 19956 16348
rect 19892 16288 19956 16292
rect 19972 16348 20036 16352
rect 19972 16292 19976 16348
rect 19976 16292 20032 16348
rect 20032 16292 20036 16348
rect 19972 16288 20036 16292
rect 23652 16348 23716 16352
rect 23652 16292 23656 16348
rect 23656 16292 23712 16348
rect 23712 16292 23716 16348
rect 23652 16288 23716 16292
rect 23732 16348 23796 16352
rect 23732 16292 23736 16348
rect 23736 16292 23792 16348
rect 23792 16292 23796 16348
rect 23732 16288 23796 16292
rect 23812 16348 23876 16352
rect 23812 16292 23816 16348
rect 23816 16292 23872 16348
rect 23872 16292 23876 16348
rect 23812 16288 23876 16292
rect 23892 16348 23956 16352
rect 23892 16292 23896 16348
rect 23896 16292 23952 16348
rect 23952 16292 23956 16348
rect 23892 16288 23956 16292
rect 23972 16348 24036 16352
rect 23972 16292 23976 16348
rect 23976 16292 24032 16348
rect 24032 16292 24036 16348
rect 23972 16288 24036 16292
rect 18644 16220 18708 16284
rect 19380 16280 19444 16284
rect 19380 16224 19394 16280
rect 19394 16224 19444 16280
rect 19380 16220 19444 16224
rect 14596 16084 14660 16148
rect 2912 15804 2976 15808
rect 2912 15748 2916 15804
rect 2916 15748 2972 15804
rect 2972 15748 2976 15804
rect 2912 15744 2976 15748
rect 2992 15804 3056 15808
rect 2992 15748 2996 15804
rect 2996 15748 3052 15804
rect 3052 15748 3056 15804
rect 2992 15744 3056 15748
rect 3072 15804 3136 15808
rect 3072 15748 3076 15804
rect 3076 15748 3132 15804
rect 3132 15748 3136 15804
rect 3072 15744 3136 15748
rect 3152 15804 3216 15808
rect 3152 15748 3156 15804
rect 3156 15748 3212 15804
rect 3212 15748 3216 15804
rect 3152 15744 3216 15748
rect 3232 15804 3296 15808
rect 3232 15748 3236 15804
rect 3236 15748 3292 15804
rect 3292 15748 3296 15804
rect 3232 15744 3296 15748
rect 6912 15804 6976 15808
rect 6912 15748 6916 15804
rect 6916 15748 6972 15804
rect 6972 15748 6976 15804
rect 6912 15744 6976 15748
rect 6992 15804 7056 15808
rect 6992 15748 6996 15804
rect 6996 15748 7052 15804
rect 7052 15748 7056 15804
rect 6992 15744 7056 15748
rect 7072 15804 7136 15808
rect 7072 15748 7076 15804
rect 7076 15748 7132 15804
rect 7132 15748 7136 15804
rect 7072 15744 7136 15748
rect 7152 15804 7216 15808
rect 7152 15748 7156 15804
rect 7156 15748 7212 15804
rect 7212 15748 7216 15804
rect 7152 15744 7216 15748
rect 7232 15804 7296 15808
rect 7232 15748 7236 15804
rect 7236 15748 7292 15804
rect 7292 15748 7296 15804
rect 7232 15744 7296 15748
rect 10912 15804 10976 15808
rect 10912 15748 10916 15804
rect 10916 15748 10972 15804
rect 10972 15748 10976 15804
rect 10912 15744 10976 15748
rect 10992 15804 11056 15808
rect 10992 15748 10996 15804
rect 10996 15748 11052 15804
rect 11052 15748 11056 15804
rect 10992 15744 11056 15748
rect 11072 15804 11136 15808
rect 11072 15748 11076 15804
rect 11076 15748 11132 15804
rect 11132 15748 11136 15804
rect 11072 15744 11136 15748
rect 11152 15804 11216 15808
rect 11152 15748 11156 15804
rect 11156 15748 11212 15804
rect 11212 15748 11216 15804
rect 11152 15744 11216 15748
rect 11232 15804 11296 15808
rect 11232 15748 11236 15804
rect 11236 15748 11292 15804
rect 11292 15748 11296 15804
rect 11232 15744 11296 15748
rect 14912 15804 14976 15808
rect 14912 15748 14916 15804
rect 14916 15748 14972 15804
rect 14972 15748 14976 15804
rect 14912 15744 14976 15748
rect 14992 15804 15056 15808
rect 14992 15748 14996 15804
rect 14996 15748 15052 15804
rect 15052 15748 15056 15804
rect 14992 15744 15056 15748
rect 15072 15804 15136 15808
rect 15072 15748 15076 15804
rect 15076 15748 15132 15804
rect 15132 15748 15136 15804
rect 15072 15744 15136 15748
rect 15152 15804 15216 15808
rect 15152 15748 15156 15804
rect 15156 15748 15212 15804
rect 15212 15748 15216 15804
rect 15152 15744 15216 15748
rect 15232 15804 15296 15808
rect 15232 15748 15236 15804
rect 15236 15748 15292 15804
rect 15292 15748 15296 15804
rect 15232 15744 15296 15748
rect 18912 15804 18976 15808
rect 18912 15748 18916 15804
rect 18916 15748 18972 15804
rect 18972 15748 18976 15804
rect 18912 15744 18976 15748
rect 18992 15804 19056 15808
rect 18992 15748 18996 15804
rect 18996 15748 19052 15804
rect 19052 15748 19056 15804
rect 18992 15744 19056 15748
rect 19072 15804 19136 15808
rect 19072 15748 19076 15804
rect 19076 15748 19132 15804
rect 19132 15748 19136 15804
rect 19072 15744 19136 15748
rect 19152 15804 19216 15808
rect 19152 15748 19156 15804
rect 19156 15748 19212 15804
rect 19212 15748 19216 15804
rect 19152 15744 19216 15748
rect 19232 15804 19296 15808
rect 19232 15748 19236 15804
rect 19236 15748 19292 15804
rect 19292 15748 19296 15804
rect 19232 15744 19296 15748
rect 22912 15804 22976 15808
rect 22912 15748 22916 15804
rect 22916 15748 22972 15804
rect 22972 15748 22976 15804
rect 22912 15744 22976 15748
rect 22992 15804 23056 15808
rect 22992 15748 22996 15804
rect 22996 15748 23052 15804
rect 23052 15748 23056 15804
rect 22992 15744 23056 15748
rect 23072 15804 23136 15808
rect 23072 15748 23076 15804
rect 23076 15748 23132 15804
rect 23132 15748 23136 15804
rect 23072 15744 23136 15748
rect 23152 15804 23216 15808
rect 23152 15748 23156 15804
rect 23156 15748 23212 15804
rect 23212 15748 23216 15804
rect 23152 15744 23216 15748
rect 23232 15804 23296 15808
rect 23232 15748 23236 15804
rect 23236 15748 23292 15804
rect 23292 15748 23296 15804
rect 23232 15744 23296 15748
rect 3652 15260 3716 15264
rect 3652 15204 3656 15260
rect 3656 15204 3712 15260
rect 3712 15204 3716 15260
rect 3652 15200 3716 15204
rect 3732 15260 3796 15264
rect 3732 15204 3736 15260
rect 3736 15204 3792 15260
rect 3792 15204 3796 15260
rect 3732 15200 3796 15204
rect 3812 15260 3876 15264
rect 3812 15204 3816 15260
rect 3816 15204 3872 15260
rect 3872 15204 3876 15260
rect 3812 15200 3876 15204
rect 3892 15260 3956 15264
rect 3892 15204 3896 15260
rect 3896 15204 3952 15260
rect 3952 15204 3956 15260
rect 3892 15200 3956 15204
rect 3972 15260 4036 15264
rect 3972 15204 3976 15260
rect 3976 15204 4032 15260
rect 4032 15204 4036 15260
rect 3972 15200 4036 15204
rect 7652 15260 7716 15264
rect 7652 15204 7656 15260
rect 7656 15204 7712 15260
rect 7712 15204 7716 15260
rect 7652 15200 7716 15204
rect 7732 15260 7796 15264
rect 7732 15204 7736 15260
rect 7736 15204 7792 15260
rect 7792 15204 7796 15260
rect 7732 15200 7796 15204
rect 7812 15260 7876 15264
rect 7812 15204 7816 15260
rect 7816 15204 7872 15260
rect 7872 15204 7876 15260
rect 7812 15200 7876 15204
rect 7892 15260 7956 15264
rect 7892 15204 7896 15260
rect 7896 15204 7952 15260
rect 7952 15204 7956 15260
rect 7892 15200 7956 15204
rect 7972 15260 8036 15264
rect 7972 15204 7976 15260
rect 7976 15204 8032 15260
rect 8032 15204 8036 15260
rect 7972 15200 8036 15204
rect 11652 15260 11716 15264
rect 11652 15204 11656 15260
rect 11656 15204 11712 15260
rect 11712 15204 11716 15260
rect 11652 15200 11716 15204
rect 11732 15260 11796 15264
rect 11732 15204 11736 15260
rect 11736 15204 11792 15260
rect 11792 15204 11796 15260
rect 11732 15200 11796 15204
rect 11812 15260 11876 15264
rect 11812 15204 11816 15260
rect 11816 15204 11872 15260
rect 11872 15204 11876 15260
rect 11812 15200 11876 15204
rect 11892 15260 11956 15264
rect 11892 15204 11896 15260
rect 11896 15204 11952 15260
rect 11952 15204 11956 15260
rect 11892 15200 11956 15204
rect 11972 15260 12036 15264
rect 11972 15204 11976 15260
rect 11976 15204 12032 15260
rect 12032 15204 12036 15260
rect 11972 15200 12036 15204
rect 15652 15260 15716 15264
rect 15652 15204 15656 15260
rect 15656 15204 15712 15260
rect 15712 15204 15716 15260
rect 15652 15200 15716 15204
rect 15732 15260 15796 15264
rect 15732 15204 15736 15260
rect 15736 15204 15792 15260
rect 15792 15204 15796 15260
rect 15732 15200 15796 15204
rect 15812 15260 15876 15264
rect 15812 15204 15816 15260
rect 15816 15204 15872 15260
rect 15872 15204 15876 15260
rect 15812 15200 15876 15204
rect 15892 15260 15956 15264
rect 15892 15204 15896 15260
rect 15896 15204 15952 15260
rect 15952 15204 15956 15260
rect 15892 15200 15956 15204
rect 15972 15260 16036 15264
rect 15972 15204 15976 15260
rect 15976 15204 16032 15260
rect 16032 15204 16036 15260
rect 15972 15200 16036 15204
rect 19652 15260 19716 15264
rect 19652 15204 19656 15260
rect 19656 15204 19712 15260
rect 19712 15204 19716 15260
rect 19652 15200 19716 15204
rect 19732 15260 19796 15264
rect 19732 15204 19736 15260
rect 19736 15204 19792 15260
rect 19792 15204 19796 15260
rect 19732 15200 19796 15204
rect 19812 15260 19876 15264
rect 19812 15204 19816 15260
rect 19816 15204 19872 15260
rect 19872 15204 19876 15260
rect 19812 15200 19876 15204
rect 19892 15260 19956 15264
rect 19892 15204 19896 15260
rect 19896 15204 19952 15260
rect 19952 15204 19956 15260
rect 19892 15200 19956 15204
rect 19972 15260 20036 15264
rect 19972 15204 19976 15260
rect 19976 15204 20032 15260
rect 20032 15204 20036 15260
rect 19972 15200 20036 15204
rect 23652 15260 23716 15264
rect 23652 15204 23656 15260
rect 23656 15204 23712 15260
rect 23712 15204 23716 15260
rect 23652 15200 23716 15204
rect 23732 15260 23796 15264
rect 23732 15204 23736 15260
rect 23736 15204 23792 15260
rect 23792 15204 23796 15260
rect 23732 15200 23796 15204
rect 23812 15260 23876 15264
rect 23812 15204 23816 15260
rect 23816 15204 23872 15260
rect 23872 15204 23876 15260
rect 23812 15200 23876 15204
rect 23892 15260 23956 15264
rect 23892 15204 23896 15260
rect 23896 15204 23952 15260
rect 23952 15204 23956 15260
rect 23892 15200 23956 15204
rect 23972 15260 24036 15264
rect 23972 15204 23976 15260
rect 23976 15204 24032 15260
rect 24032 15204 24036 15260
rect 23972 15200 24036 15204
rect 2912 14716 2976 14720
rect 2912 14660 2916 14716
rect 2916 14660 2972 14716
rect 2972 14660 2976 14716
rect 2912 14656 2976 14660
rect 2992 14716 3056 14720
rect 2992 14660 2996 14716
rect 2996 14660 3052 14716
rect 3052 14660 3056 14716
rect 2992 14656 3056 14660
rect 3072 14716 3136 14720
rect 3072 14660 3076 14716
rect 3076 14660 3132 14716
rect 3132 14660 3136 14716
rect 3072 14656 3136 14660
rect 3152 14716 3216 14720
rect 3152 14660 3156 14716
rect 3156 14660 3212 14716
rect 3212 14660 3216 14716
rect 3152 14656 3216 14660
rect 3232 14716 3296 14720
rect 3232 14660 3236 14716
rect 3236 14660 3292 14716
rect 3292 14660 3296 14716
rect 3232 14656 3296 14660
rect 6912 14716 6976 14720
rect 6912 14660 6916 14716
rect 6916 14660 6972 14716
rect 6972 14660 6976 14716
rect 6912 14656 6976 14660
rect 6992 14716 7056 14720
rect 6992 14660 6996 14716
rect 6996 14660 7052 14716
rect 7052 14660 7056 14716
rect 6992 14656 7056 14660
rect 7072 14716 7136 14720
rect 7072 14660 7076 14716
rect 7076 14660 7132 14716
rect 7132 14660 7136 14716
rect 7072 14656 7136 14660
rect 7152 14716 7216 14720
rect 7152 14660 7156 14716
rect 7156 14660 7212 14716
rect 7212 14660 7216 14716
rect 7152 14656 7216 14660
rect 7232 14716 7296 14720
rect 7232 14660 7236 14716
rect 7236 14660 7292 14716
rect 7292 14660 7296 14716
rect 7232 14656 7296 14660
rect 10912 14716 10976 14720
rect 10912 14660 10916 14716
rect 10916 14660 10972 14716
rect 10972 14660 10976 14716
rect 10912 14656 10976 14660
rect 10992 14716 11056 14720
rect 10992 14660 10996 14716
rect 10996 14660 11052 14716
rect 11052 14660 11056 14716
rect 10992 14656 11056 14660
rect 11072 14716 11136 14720
rect 11072 14660 11076 14716
rect 11076 14660 11132 14716
rect 11132 14660 11136 14716
rect 11072 14656 11136 14660
rect 11152 14716 11216 14720
rect 11152 14660 11156 14716
rect 11156 14660 11212 14716
rect 11212 14660 11216 14716
rect 11152 14656 11216 14660
rect 11232 14716 11296 14720
rect 11232 14660 11236 14716
rect 11236 14660 11292 14716
rect 11292 14660 11296 14716
rect 11232 14656 11296 14660
rect 14912 14716 14976 14720
rect 14912 14660 14916 14716
rect 14916 14660 14972 14716
rect 14972 14660 14976 14716
rect 14912 14656 14976 14660
rect 14992 14716 15056 14720
rect 14992 14660 14996 14716
rect 14996 14660 15052 14716
rect 15052 14660 15056 14716
rect 14992 14656 15056 14660
rect 15072 14716 15136 14720
rect 15072 14660 15076 14716
rect 15076 14660 15132 14716
rect 15132 14660 15136 14716
rect 15072 14656 15136 14660
rect 15152 14716 15216 14720
rect 15152 14660 15156 14716
rect 15156 14660 15212 14716
rect 15212 14660 15216 14716
rect 15152 14656 15216 14660
rect 15232 14716 15296 14720
rect 15232 14660 15236 14716
rect 15236 14660 15292 14716
rect 15292 14660 15296 14716
rect 15232 14656 15296 14660
rect 18912 14716 18976 14720
rect 18912 14660 18916 14716
rect 18916 14660 18972 14716
rect 18972 14660 18976 14716
rect 18912 14656 18976 14660
rect 18992 14716 19056 14720
rect 18992 14660 18996 14716
rect 18996 14660 19052 14716
rect 19052 14660 19056 14716
rect 18992 14656 19056 14660
rect 19072 14716 19136 14720
rect 19072 14660 19076 14716
rect 19076 14660 19132 14716
rect 19132 14660 19136 14716
rect 19072 14656 19136 14660
rect 19152 14716 19216 14720
rect 19152 14660 19156 14716
rect 19156 14660 19212 14716
rect 19212 14660 19216 14716
rect 19152 14656 19216 14660
rect 19232 14716 19296 14720
rect 19232 14660 19236 14716
rect 19236 14660 19292 14716
rect 19292 14660 19296 14716
rect 19232 14656 19296 14660
rect 22912 14716 22976 14720
rect 22912 14660 22916 14716
rect 22916 14660 22972 14716
rect 22972 14660 22976 14716
rect 22912 14656 22976 14660
rect 22992 14716 23056 14720
rect 22992 14660 22996 14716
rect 22996 14660 23052 14716
rect 23052 14660 23056 14716
rect 22992 14656 23056 14660
rect 23072 14716 23136 14720
rect 23072 14660 23076 14716
rect 23076 14660 23132 14716
rect 23132 14660 23136 14716
rect 23072 14656 23136 14660
rect 23152 14716 23216 14720
rect 23152 14660 23156 14716
rect 23156 14660 23212 14716
rect 23212 14660 23216 14716
rect 23152 14656 23216 14660
rect 23232 14716 23296 14720
rect 23232 14660 23236 14716
rect 23236 14660 23292 14716
rect 23292 14660 23296 14716
rect 23232 14656 23296 14660
rect 14596 14452 14660 14516
rect 15516 14452 15580 14516
rect 18276 14316 18340 14380
rect 3652 14172 3716 14176
rect 3652 14116 3656 14172
rect 3656 14116 3712 14172
rect 3712 14116 3716 14172
rect 3652 14112 3716 14116
rect 3732 14172 3796 14176
rect 3732 14116 3736 14172
rect 3736 14116 3792 14172
rect 3792 14116 3796 14172
rect 3732 14112 3796 14116
rect 3812 14172 3876 14176
rect 3812 14116 3816 14172
rect 3816 14116 3872 14172
rect 3872 14116 3876 14172
rect 3812 14112 3876 14116
rect 3892 14172 3956 14176
rect 3892 14116 3896 14172
rect 3896 14116 3952 14172
rect 3952 14116 3956 14172
rect 3892 14112 3956 14116
rect 3972 14172 4036 14176
rect 3972 14116 3976 14172
rect 3976 14116 4032 14172
rect 4032 14116 4036 14172
rect 3972 14112 4036 14116
rect 7652 14172 7716 14176
rect 7652 14116 7656 14172
rect 7656 14116 7712 14172
rect 7712 14116 7716 14172
rect 7652 14112 7716 14116
rect 7732 14172 7796 14176
rect 7732 14116 7736 14172
rect 7736 14116 7792 14172
rect 7792 14116 7796 14172
rect 7732 14112 7796 14116
rect 7812 14172 7876 14176
rect 7812 14116 7816 14172
rect 7816 14116 7872 14172
rect 7872 14116 7876 14172
rect 7812 14112 7876 14116
rect 7892 14172 7956 14176
rect 7892 14116 7896 14172
rect 7896 14116 7952 14172
rect 7952 14116 7956 14172
rect 7892 14112 7956 14116
rect 7972 14172 8036 14176
rect 7972 14116 7976 14172
rect 7976 14116 8032 14172
rect 8032 14116 8036 14172
rect 7972 14112 8036 14116
rect 11652 14172 11716 14176
rect 11652 14116 11656 14172
rect 11656 14116 11712 14172
rect 11712 14116 11716 14172
rect 11652 14112 11716 14116
rect 11732 14172 11796 14176
rect 11732 14116 11736 14172
rect 11736 14116 11792 14172
rect 11792 14116 11796 14172
rect 11732 14112 11796 14116
rect 11812 14172 11876 14176
rect 11812 14116 11816 14172
rect 11816 14116 11872 14172
rect 11872 14116 11876 14172
rect 11812 14112 11876 14116
rect 11892 14172 11956 14176
rect 11892 14116 11896 14172
rect 11896 14116 11952 14172
rect 11952 14116 11956 14172
rect 11892 14112 11956 14116
rect 11972 14172 12036 14176
rect 11972 14116 11976 14172
rect 11976 14116 12032 14172
rect 12032 14116 12036 14172
rect 11972 14112 12036 14116
rect 15652 14172 15716 14176
rect 15652 14116 15656 14172
rect 15656 14116 15712 14172
rect 15712 14116 15716 14172
rect 15652 14112 15716 14116
rect 15732 14172 15796 14176
rect 15732 14116 15736 14172
rect 15736 14116 15792 14172
rect 15792 14116 15796 14172
rect 15732 14112 15796 14116
rect 15812 14172 15876 14176
rect 15812 14116 15816 14172
rect 15816 14116 15872 14172
rect 15872 14116 15876 14172
rect 15812 14112 15876 14116
rect 15892 14172 15956 14176
rect 15892 14116 15896 14172
rect 15896 14116 15952 14172
rect 15952 14116 15956 14172
rect 15892 14112 15956 14116
rect 15972 14172 16036 14176
rect 15972 14116 15976 14172
rect 15976 14116 16032 14172
rect 16032 14116 16036 14172
rect 15972 14112 16036 14116
rect 19652 14172 19716 14176
rect 19652 14116 19656 14172
rect 19656 14116 19712 14172
rect 19712 14116 19716 14172
rect 19652 14112 19716 14116
rect 19732 14172 19796 14176
rect 19732 14116 19736 14172
rect 19736 14116 19792 14172
rect 19792 14116 19796 14172
rect 19732 14112 19796 14116
rect 19812 14172 19876 14176
rect 19812 14116 19816 14172
rect 19816 14116 19872 14172
rect 19872 14116 19876 14172
rect 19812 14112 19876 14116
rect 19892 14172 19956 14176
rect 19892 14116 19896 14172
rect 19896 14116 19952 14172
rect 19952 14116 19956 14172
rect 19892 14112 19956 14116
rect 19972 14172 20036 14176
rect 19972 14116 19976 14172
rect 19976 14116 20032 14172
rect 20032 14116 20036 14172
rect 19972 14112 20036 14116
rect 23652 14172 23716 14176
rect 23652 14116 23656 14172
rect 23656 14116 23712 14172
rect 23712 14116 23716 14172
rect 23652 14112 23716 14116
rect 23732 14172 23796 14176
rect 23732 14116 23736 14172
rect 23736 14116 23792 14172
rect 23792 14116 23796 14172
rect 23732 14112 23796 14116
rect 23812 14172 23876 14176
rect 23812 14116 23816 14172
rect 23816 14116 23872 14172
rect 23872 14116 23876 14172
rect 23812 14112 23876 14116
rect 23892 14172 23956 14176
rect 23892 14116 23896 14172
rect 23896 14116 23952 14172
rect 23952 14116 23956 14172
rect 23892 14112 23956 14116
rect 23972 14172 24036 14176
rect 23972 14116 23976 14172
rect 23976 14116 24032 14172
rect 24032 14116 24036 14172
rect 23972 14112 24036 14116
rect 2912 13628 2976 13632
rect 2912 13572 2916 13628
rect 2916 13572 2972 13628
rect 2972 13572 2976 13628
rect 2912 13568 2976 13572
rect 2992 13628 3056 13632
rect 2992 13572 2996 13628
rect 2996 13572 3052 13628
rect 3052 13572 3056 13628
rect 2992 13568 3056 13572
rect 3072 13628 3136 13632
rect 3072 13572 3076 13628
rect 3076 13572 3132 13628
rect 3132 13572 3136 13628
rect 3072 13568 3136 13572
rect 3152 13628 3216 13632
rect 3152 13572 3156 13628
rect 3156 13572 3212 13628
rect 3212 13572 3216 13628
rect 3152 13568 3216 13572
rect 3232 13628 3296 13632
rect 3232 13572 3236 13628
rect 3236 13572 3292 13628
rect 3292 13572 3296 13628
rect 3232 13568 3296 13572
rect 6912 13628 6976 13632
rect 6912 13572 6916 13628
rect 6916 13572 6972 13628
rect 6972 13572 6976 13628
rect 6912 13568 6976 13572
rect 6992 13628 7056 13632
rect 6992 13572 6996 13628
rect 6996 13572 7052 13628
rect 7052 13572 7056 13628
rect 6992 13568 7056 13572
rect 7072 13628 7136 13632
rect 7072 13572 7076 13628
rect 7076 13572 7132 13628
rect 7132 13572 7136 13628
rect 7072 13568 7136 13572
rect 7152 13628 7216 13632
rect 7152 13572 7156 13628
rect 7156 13572 7212 13628
rect 7212 13572 7216 13628
rect 7152 13568 7216 13572
rect 7232 13628 7296 13632
rect 7232 13572 7236 13628
rect 7236 13572 7292 13628
rect 7292 13572 7296 13628
rect 7232 13568 7296 13572
rect 10912 13628 10976 13632
rect 10912 13572 10916 13628
rect 10916 13572 10972 13628
rect 10972 13572 10976 13628
rect 10912 13568 10976 13572
rect 10992 13628 11056 13632
rect 10992 13572 10996 13628
rect 10996 13572 11052 13628
rect 11052 13572 11056 13628
rect 10992 13568 11056 13572
rect 11072 13628 11136 13632
rect 11072 13572 11076 13628
rect 11076 13572 11132 13628
rect 11132 13572 11136 13628
rect 11072 13568 11136 13572
rect 11152 13628 11216 13632
rect 11152 13572 11156 13628
rect 11156 13572 11212 13628
rect 11212 13572 11216 13628
rect 11152 13568 11216 13572
rect 11232 13628 11296 13632
rect 11232 13572 11236 13628
rect 11236 13572 11292 13628
rect 11292 13572 11296 13628
rect 11232 13568 11296 13572
rect 14912 13628 14976 13632
rect 14912 13572 14916 13628
rect 14916 13572 14972 13628
rect 14972 13572 14976 13628
rect 14912 13568 14976 13572
rect 14992 13628 15056 13632
rect 14992 13572 14996 13628
rect 14996 13572 15052 13628
rect 15052 13572 15056 13628
rect 14992 13568 15056 13572
rect 15072 13628 15136 13632
rect 15072 13572 15076 13628
rect 15076 13572 15132 13628
rect 15132 13572 15136 13628
rect 15072 13568 15136 13572
rect 15152 13628 15216 13632
rect 15152 13572 15156 13628
rect 15156 13572 15212 13628
rect 15212 13572 15216 13628
rect 15152 13568 15216 13572
rect 15232 13628 15296 13632
rect 15232 13572 15236 13628
rect 15236 13572 15292 13628
rect 15292 13572 15296 13628
rect 15232 13568 15296 13572
rect 18912 13628 18976 13632
rect 18912 13572 18916 13628
rect 18916 13572 18972 13628
rect 18972 13572 18976 13628
rect 18912 13568 18976 13572
rect 18992 13628 19056 13632
rect 18992 13572 18996 13628
rect 18996 13572 19052 13628
rect 19052 13572 19056 13628
rect 18992 13568 19056 13572
rect 19072 13628 19136 13632
rect 19072 13572 19076 13628
rect 19076 13572 19132 13628
rect 19132 13572 19136 13628
rect 19072 13568 19136 13572
rect 19152 13628 19216 13632
rect 19152 13572 19156 13628
rect 19156 13572 19212 13628
rect 19212 13572 19216 13628
rect 19152 13568 19216 13572
rect 19232 13628 19296 13632
rect 19232 13572 19236 13628
rect 19236 13572 19292 13628
rect 19292 13572 19296 13628
rect 19232 13568 19296 13572
rect 22912 13628 22976 13632
rect 22912 13572 22916 13628
rect 22916 13572 22972 13628
rect 22972 13572 22976 13628
rect 22912 13568 22976 13572
rect 22992 13628 23056 13632
rect 22992 13572 22996 13628
rect 22996 13572 23052 13628
rect 23052 13572 23056 13628
rect 22992 13568 23056 13572
rect 23072 13628 23136 13632
rect 23072 13572 23076 13628
rect 23076 13572 23132 13628
rect 23132 13572 23136 13628
rect 23072 13568 23136 13572
rect 23152 13628 23216 13632
rect 23152 13572 23156 13628
rect 23156 13572 23212 13628
rect 23212 13572 23216 13628
rect 23152 13568 23216 13572
rect 23232 13628 23296 13632
rect 23232 13572 23236 13628
rect 23236 13572 23292 13628
rect 23292 13572 23296 13628
rect 23232 13568 23296 13572
rect 18460 13424 18524 13428
rect 18460 13368 18474 13424
rect 18474 13368 18524 13424
rect 18460 13364 18524 13368
rect 3652 13084 3716 13088
rect 3652 13028 3656 13084
rect 3656 13028 3712 13084
rect 3712 13028 3716 13084
rect 3652 13024 3716 13028
rect 3732 13084 3796 13088
rect 3732 13028 3736 13084
rect 3736 13028 3792 13084
rect 3792 13028 3796 13084
rect 3732 13024 3796 13028
rect 3812 13084 3876 13088
rect 3812 13028 3816 13084
rect 3816 13028 3872 13084
rect 3872 13028 3876 13084
rect 3812 13024 3876 13028
rect 3892 13084 3956 13088
rect 3892 13028 3896 13084
rect 3896 13028 3952 13084
rect 3952 13028 3956 13084
rect 3892 13024 3956 13028
rect 3972 13084 4036 13088
rect 3972 13028 3976 13084
rect 3976 13028 4032 13084
rect 4032 13028 4036 13084
rect 3972 13024 4036 13028
rect 7652 13084 7716 13088
rect 7652 13028 7656 13084
rect 7656 13028 7712 13084
rect 7712 13028 7716 13084
rect 7652 13024 7716 13028
rect 7732 13084 7796 13088
rect 7732 13028 7736 13084
rect 7736 13028 7792 13084
rect 7792 13028 7796 13084
rect 7732 13024 7796 13028
rect 7812 13084 7876 13088
rect 7812 13028 7816 13084
rect 7816 13028 7872 13084
rect 7872 13028 7876 13084
rect 7812 13024 7876 13028
rect 7892 13084 7956 13088
rect 7892 13028 7896 13084
rect 7896 13028 7952 13084
rect 7952 13028 7956 13084
rect 7892 13024 7956 13028
rect 7972 13084 8036 13088
rect 7972 13028 7976 13084
rect 7976 13028 8032 13084
rect 8032 13028 8036 13084
rect 7972 13024 8036 13028
rect 11652 13084 11716 13088
rect 11652 13028 11656 13084
rect 11656 13028 11712 13084
rect 11712 13028 11716 13084
rect 11652 13024 11716 13028
rect 11732 13084 11796 13088
rect 11732 13028 11736 13084
rect 11736 13028 11792 13084
rect 11792 13028 11796 13084
rect 11732 13024 11796 13028
rect 11812 13084 11876 13088
rect 11812 13028 11816 13084
rect 11816 13028 11872 13084
rect 11872 13028 11876 13084
rect 11812 13024 11876 13028
rect 11892 13084 11956 13088
rect 11892 13028 11896 13084
rect 11896 13028 11952 13084
rect 11952 13028 11956 13084
rect 11892 13024 11956 13028
rect 11972 13084 12036 13088
rect 11972 13028 11976 13084
rect 11976 13028 12032 13084
rect 12032 13028 12036 13084
rect 11972 13024 12036 13028
rect 15652 13084 15716 13088
rect 15652 13028 15656 13084
rect 15656 13028 15712 13084
rect 15712 13028 15716 13084
rect 15652 13024 15716 13028
rect 15732 13084 15796 13088
rect 15732 13028 15736 13084
rect 15736 13028 15792 13084
rect 15792 13028 15796 13084
rect 15732 13024 15796 13028
rect 15812 13084 15876 13088
rect 15812 13028 15816 13084
rect 15816 13028 15872 13084
rect 15872 13028 15876 13084
rect 15812 13024 15876 13028
rect 15892 13084 15956 13088
rect 15892 13028 15896 13084
rect 15896 13028 15952 13084
rect 15952 13028 15956 13084
rect 15892 13024 15956 13028
rect 15972 13084 16036 13088
rect 15972 13028 15976 13084
rect 15976 13028 16032 13084
rect 16032 13028 16036 13084
rect 15972 13024 16036 13028
rect 19652 13084 19716 13088
rect 19652 13028 19656 13084
rect 19656 13028 19712 13084
rect 19712 13028 19716 13084
rect 19652 13024 19716 13028
rect 19732 13084 19796 13088
rect 19732 13028 19736 13084
rect 19736 13028 19792 13084
rect 19792 13028 19796 13084
rect 19732 13024 19796 13028
rect 19812 13084 19876 13088
rect 19812 13028 19816 13084
rect 19816 13028 19872 13084
rect 19872 13028 19876 13084
rect 19812 13024 19876 13028
rect 19892 13084 19956 13088
rect 19892 13028 19896 13084
rect 19896 13028 19952 13084
rect 19952 13028 19956 13084
rect 19892 13024 19956 13028
rect 19972 13084 20036 13088
rect 19972 13028 19976 13084
rect 19976 13028 20032 13084
rect 20032 13028 20036 13084
rect 19972 13024 20036 13028
rect 23652 13084 23716 13088
rect 23652 13028 23656 13084
rect 23656 13028 23712 13084
rect 23712 13028 23716 13084
rect 23652 13024 23716 13028
rect 23732 13084 23796 13088
rect 23732 13028 23736 13084
rect 23736 13028 23792 13084
rect 23792 13028 23796 13084
rect 23732 13024 23796 13028
rect 23812 13084 23876 13088
rect 23812 13028 23816 13084
rect 23816 13028 23872 13084
rect 23872 13028 23876 13084
rect 23812 13024 23876 13028
rect 23892 13084 23956 13088
rect 23892 13028 23896 13084
rect 23896 13028 23952 13084
rect 23952 13028 23956 13084
rect 23892 13024 23956 13028
rect 23972 13084 24036 13088
rect 23972 13028 23976 13084
rect 23976 13028 24032 13084
rect 24032 13028 24036 13084
rect 23972 13024 24036 13028
rect 5212 12880 5276 12884
rect 5212 12824 5262 12880
rect 5262 12824 5276 12880
rect 5212 12820 5276 12824
rect 2912 12540 2976 12544
rect 2912 12484 2916 12540
rect 2916 12484 2972 12540
rect 2972 12484 2976 12540
rect 2912 12480 2976 12484
rect 2992 12540 3056 12544
rect 2992 12484 2996 12540
rect 2996 12484 3052 12540
rect 3052 12484 3056 12540
rect 2992 12480 3056 12484
rect 3072 12540 3136 12544
rect 3072 12484 3076 12540
rect 3076 12484 3132 12540
rect 3132 12484 3136 12540
rect 3072 12480 3136 12484
rect 3152 12540 3216 12544
rect 3152 12484 3156 12540
rect 3156 12484 3212 12540
rect 3212 12484 3216 12540
rect 3152 12480 3216 12484
rect 3232 12540 3296 12544
rect 3232 12484 3236 12540
rect 3236 12484 3292 12540
rect 3292 12484 3296 12540
rect 3232 12480 3296 12484
rect 6912 12540 6976 12544
rect 6912 12484 6916 12540
rect 6916 12484 6972 12540
rect 6972 12484 6976 12540
rect 6912 12480 6976 12484
rect 6992 12540 7056 12544
rect 6992 12484 6996 12540
rect 6996 12484 7052 12540
rect 7052 12484 7056 12540
rect 6992 12480 7056 12484
rect 7072 12540 7136 12544
rect 7072 12484 7076 12540
rect 7076 12484 7132 12540
rect 7132 12484 7136 12540
rect 7072 12480 7136 12484
rect 7152 12540 7216 12544
rect 7152 12484 7156 12540
rect 7156 12484 7212 12540
rect 7212 12484 7216 12540
rect 7152 12480 7216 12484
rect 7232 12540 7296 12544
rect 7232 12484 7236 12540
rect 7236 12484 7292 12540
rect 7292 12484 7296 12540
rect 7232 12480 7296 12484
rect 10912 12540 10976 12544
rect 10912 12484 10916 12540
rect 10916 12484 10972 12540
rect 10972 12484 10976 12540
rect 10912 12480 10976 12484
rect 10992 12540 11056 12544
rect 10992 12484 10996 12540
rect 10996 12484 11052 12540
rect 11052 12484 11056 12540
rect 10992 12480 11056 12484
rect 11072 12540 11136 12544
rect 11072 12484 11076 12540
rect 11076 12484 11132 12540
rect 11132 12484 11136 12540
rect 11072 12480 11136 12484
rect 11152 12540 11216 12544
rect 11152 12484 11156 12540
rect 11156 12484 11212 12540
rect 11212 12484 11216 12540
rect 11152 12480 11216 12484
rect 11232 12540 11296 12544
rect 11232 12484 11236 12540
rect 11236 12484 11292 12540
rect 11292 12484 11296 12540
rect 11232 12480 11296 12484
rect 14912 12540 14976 12544
rect 14912 12484 14916 12540
rect 14916 12484 14972 12540
rect 14972 12484 14976 12540
rect 14912 12480 14976 12484
rect 14992 12540 15056 12544
rect 14992 12484 14996 12540
rect 14996 12484 15052 12540
rect 15052 12484 15056 12540
rect 14992 12480 15056 12484
rect 15072 12540 15136 12544
rect 15072 12484 15076 12540
rect 15076 12484 15132 12540
rect 15132 12484 15136 12540
rect 15072 12480 15136 12484
rect 15152 12540 15216 12544
rect 15152 12484 15156 12540
rect 15156 12484 15212 12540
rect 15212 12484 15216 12540
rect 15152 12480 15216 12484
rect 15232 12540 15296 12544
rect 15232 12484 15236 12540
rect 15236 12484 15292 12540
rect 15292 12484 15296 12540
rect 15232 12480 15296 12484
rect 18912 12540 18976 12544
rect 18912 12484 18916 12540
rect 18916 12484 18972 12540
rect 18972 12484 18976 12540
rect 18912 12480 18976 12484
rect 18992 12540 19056 12544
rect 18992 12484 18996 12540
rect 18996 12484 19052 12540
rect 19052 12484 19056 12540
rect 18992 12480 19056 12484
rect 19072 12540 19136 12544
rect 19072 12484 19076 12540
rect 19076 12484 19132 12540
rect 19132 12484 19136 12540
rect 19072 12480 19136 12484
rect 19152 12540 19216 12544
rect 19152 12484 19156 12540
rect 19156 12484 19212 12540
rect 19212 12484 19216 12540
rect 19152 12480 19216 12484
rect 19232 12540 19296 12544
rect 19232 12484 19236 12540
rect 19236 12484 19292 12540
rect 19292 12484 19296 12540
rect 19232 12480 19296 12484
rect 22912 12540 22976 12544
rect 22912 12484 22916 12540
rect 22916 12484 22972 12540
rect 22972 12484 22976 12540
rect 22912 12480 22976 12484
rect 22992 12540 23056 12544
rect 22992 12484 22996 12540
rect 22996 12484 23052 12540
rect 23052 12484 23056 12540
rect 22992 12480 23056 12484
rect 23072 12540 23136 12544
rect 23072 12484 23076 12540
rect 23076 12484 23132 12540
rect 23132 12484 23136 12540
rect 23072 12480 23136 12484
rect 23152 12540 23216 12544
rect 23152 12484 23156 12540
rect 23156 12484 23212 12540
rect 23212 12484 23216 12540
rect 23152 12480 23216 12484
rect 23232 12540 23296 12544
rect 23232 12484 23236 12540
rect 23236 12484 23292 12540
rect 23292 12484 23296 12540
rect 23232 12480 23296 12484
rect 3652 11996 3716 12000
rect 3652 11940 3656 11996
rect 3656 11940 3712 11996
rect 3712 11940 3716 11996
rect 3652 11936 3716 11940
rect 3732 11996 3796 12000
rect 3732 11940 3736 11996
rect 3736 11940 3792 11996
rect 3792 11940 3796 11996
rect 3732 11936 3796 11940
rect 3812 11996 3876 12000
rect 3812 11940 3816 11996
rect 3816 11940 3872 11996
rect 3872 11940 3876 11996
rect 3812 11936 3876 11940
rect 3892 11996 3956 12000
rect 3892 11940 3896 11996
rect 3896 11940 3952 11996
rect 3952 11940 3956 11996
rect 3892 11936 3956 11940
rect 3972 11996 4036 12000
rect 3972 11940 3976 11996
rect 3976 11940 4032 11996
rect 4032 11940 4036 11996
rect 3972 11936 4036 11940
rect 7652 11996 7716 12000
rect 7652 11940 7656 11996
rect 7656 11940 7712 11996
rect 7712 11940 7716 11996
rect 7652 11936 7716 11940
rect 7732 11996 7796 12000
rect 7732 11940 7736 11996
rect 7736 11940 7792 11996
rect 7792 11940 7796 11996
rect 7732 11936 7796 11940
rect 7812 11996 7876 12000
rect 7812 11940 7816 11996
rect 7816 11940 7872 11996
rect 7872 11940 7876 11996
rect 7812 11936 7876 11940
rect 7892 11996 7956 12000
rect 7892 11940 7896 11996
rect 7896 11940 7952 11996
rect 7952 11940 7956 11996
rect 7892 11936 7956 11940
rect 7972 11996 8036 12000
rect 7972 11940 7976 11996
rect 7976 11940 8032 11996
rect 8032 11940 8036 11996
rect 7972 11936 8036 11940
rect 11652 11996 11716 12000
rect 11652 11940 11656 11996
rect 11656 11940 11712 11996
rect 11712 11940 11716 11996
rect 11652 11936 11716 11940
rect 11732 11996 11796 12000
rect 11732 11940 11736 11996
rect 11736 11940 11792 11996
rect 11792 11940 11796 11996
rect 11732 11936 11796 11940
rect 11812 11996 11876 12000
rect 11812 11940 11816 11996
rect 11816 11940 11872 11996
rect 11872 11940 11876 11996
rect 11812 11936 11876 11940
rect 11892 11996 11956 12000
rect 11892 11940 11896 11996
rect 11896 11940 11952 11996
rect 11952 11940 11956 11996
rect 11892 11936 11956 11940
rect 11972 11996 12036 12000
rect 11972 11940 11976 11996
rect 11976 11940 12032 11996
rect 12032 11940 12036 11996
rect 11972 11936 12036 11940
rect 15652 11996 15716 12000
rect 15652 11940 15656 11996
rect 15656 11940 15712 11996
rect 15712 11940 15716 11996
rect 15652 11936 15716 11940
rect 15732 11996 15796 12000
rect 15732 11940 15736 11996
rect 15736 11940 15792 11996
rect 15792 11940 15796 11996
rect 15732 11936 15796 11940
rect 15812 11996 15876 12000
rect 15812 11940 15816 11996
rect 15816 11940 15872 11996
rect 15872 11940 15876 11996
rect 15812 11936 15876 11940
rect 15892 11996 15956 12000
rect 15892 11940 15896 11996
rect 15896 11940 15952 11996
rect 15952 11940 15956 11996
rect 15892 11936 15956 11940
rect 15972 11996 16036 12000
rect 15972 11940 15976 11996
rect 15976 11940 16032 11996
rect 16032 11940 16036 11996
rect 15972 11936 16036 11940
rect 19652 11996 19716 12000
rect 19652 11940 19656 11996
rect 19656 11940 19712 11996
rect 19712 11940 19716 11996
rect 19652 11936 19716 11940
rect 19732 11996 19796 12000
rect 19732 11940 19736 11996
rect 19736 11940 19792 11996
rect 19792 11940 19796 11996
rect 19732 11936 19796 11940
rect 19812 11996 19876 12000
rect 19812 11940 19816 11996
rect 19816 11940 19872 11996
rect 19872 11940 19876 11996
rect 19812 11936 19876 11940
rect 19892 11996 19956 12000
rect 19892 11940 19896 11996
rect 19896 11940 19952 11996
rect 19952 11940 19956 11996
rect 19892 11936 19956 11940
rect 19972 11996 20036 12000
rect 19972 11940 19976 11996
rect 19976 11940 20032 11996
rect 20032 11940 20036 11996
rect 19972 11936 20036 11940
rect 23652 11996 23716 12000
rect 23652 11940 23656 11996
rect 23656 11940 23712 11996
rect 23712 11940 23716 11996
rect 23652 11936 23716 11940
rect 23732 11996 23796 12000
rect 23732 11940 23736 11996
rect 23736 11940 23792 11996
rect 23792 11940 23796 11996
rect 23732 11936 23796 11940
rect 23812 11996 23876 12000
rect 23812 11940 23816 11996
rect 23816 11940 23872 11996
rect 23872 11940 23876 11996
rect 23812 11936 23876 11940
rect 23892 11996 23956 12000
rect 23892 11940 23896 11996
rect 23896 11940 23952 11996
rect 23952 11940 23956 11996
rect 23892 11936 23956 11940
rect 23972 11996 24036 12000
rect 23972 11940 23976 11996
rect 23976 11940 24032 11996
rect 24032 11940 24036 11996
rect 23972 11936 24036 11940
rect 5396 11732 5460 11796
rect 9996 11596 10060 11660
rect 2912 11452 2976 11456
rect 2912 11396 2916 11452
rect 2916 11396 2972 11452
rect 2972 11396 2976 11452
rect 2912 11392 2976 11396
rect 2992 11452 3056 11456
rect 2992 11396 2996 11452
rect 2996 11396 3052 11452
rect 3052 11396 3056 11452
rect 2992 11392 3056 11396
rect 3072 11452 3136 11456
rect 3072 11396 3076 11452
rect 3076 11396 3132 11452
rect 3132 11396 3136 11452
rect 3072 11392 3136 11396
rect 3152 11452 3216 11456
rect 3152 11396 3156 11452
rect 3156 11396 3212 11452
rect 3212 11396 3216 11452
rect 3152 11392 3216 11396
rect 3232 11452 3296 11456
rect 3232 11396 3236 11452
rect 3236 11396 3292 11452
rect 3292 11396 3296 11452
rect 3232 11392 3296 11396
rect 6912 11452 6976 11456
rect 6912 11396 6916 11452
rect 6916 11396 6972 11452
rect 6972 11396 6976 11452
rect 6912 11392 6976 11396
rect 6992 11452 7056 11456
rect 6992 11396 6996 11452
rect 6996 11396 7052 11452
rect 7052 11396 7056 11452
rect 6992 11392 7056 11396
rect 7072 11452 7136 11456
rect 7072 11396 7076 11452
rect 7076 11396 7132 11452
rect 7132 11396 7136 11452
rect 7072 11392 7136 11396
rect 7152 11452 7216 11456
rect 7152 11396 7156 11452
rect 7156 11396 7212 11452
rect 7212 11396 7216 11452
rect 7152 11392 7216 11396
rect 7232 11452 7296 11456
rect 7232 11396 7236 11452
rect 7236 11396 7292 11452
rect 7292 11396 7296 11452
rect 7232 11392 7296 11396
rect 10912 11452 10976 11456
rect 10912 11396 10916 11452
rect 10916 11396 10972 11452
rect 10972 11396 10976 11452
rect 10912 11392 10976 11396
rect 10992 11452 11056 11456
rect 10992 11396 10996 11452
rect 10996 11396 11052 11452
rect 11052 11396 11056 11452
rect 10992 11392 11056 11396
rect 11072 11452 11136 11456
rect 11072 11396 11076 11452
rect 11076 11396 11132 11452
rect 11132 11396 11136 11452
rect 11072 11392 11136 11396
rect 11152 11452 11216 11456
rect 11152 11396 11156 11452
rect 11156 11396 11212 11452
rect 11212 11396 11216 11452
rect 11152 11392 11216 11396
rect 11232 11452 11296 11456
rect 11232 11396 11236 11452
rect 11236 11396 11292 11452
rect 11292 11396 11296 11452
rect 11232 11392 11296 11396
rect 14912 11452 14976 11456
rect 14912 11396 14916 11452
rect 14916 11396 14972 11452
rect 14972 11396 14976 11452
rect 14912 11392 14976 11396
rect 14992 11452 15056 11456
rect 14992 11396 14996 11452
rect 14996 11396 15052 11452
rect 15052 11396 15056 11452
rect 14992 11392 15056 11396
rect 15072 11452 15136 11456
rect 15072 11396 15076 11452
rect 15076 11396 15132 11452
rect 15132 11396 15136 11452
rect 15072 11392 15136 11396
rect 15152 11452 15216 11456
rect 15152 11396 15156 11452
rect 15156 11396 15212 11452
rect 15212 11396 15216 11452
rect 15152 11392 15216 11396
rect 15232 11452 15296 11456
rect 15232 11396 15236 11452
rect 15236 11396 15292 11452
rect 15292 11396 15296 11452
rect 15232 11392 15296 11396
rect 18912 11452 18976 11456
rect 18912 11396 18916 11452
rect 18916 11396 18972 11452
rect 18972 11396 18976 11452
rect 18912 11392 18976 11396
rect 18992 11452 19056 11456
rect 18992 11396 18996 11452
rect 18996 11396 19052 11452
rect 19052 11396 19056 11452
rect 18992 11392 19056 11396
rect 19072 11452 19136 11456
rect 19072 11396 19076 11452
rect 19076 11396 19132 11452
rect 19132 11396 19136 11452
rect 19072 11392 19136 11396
rect 19152 11452 19216 11456
rect 19152 11396 19156 11452
rect 19156 11396 19212 11452
rect 19212 11396 19216 11452
rect 19152 11392 19216 11396
rect 19232 11452 19296 11456
rect 19232 11396 19236 11452
rect 19236 11396 19292 11452
rect 19292 11396 19296 11452
rect 19232 11392 19296 11396
rect 22912 11452 22976 11456
rect 22912 11396 22916 11452
rect 22916 11396 22972 11452
rect 22972 11396 22976 11452
rect 22912 11392 22976 11396
rect 22992 11452 23056 11456
rect 22992 11396 22996 11452
rect 22996 11396 23052 11452
rect 23052 11396 23056 11452
rect 22992 11392 23056 11396
rect 23072 11452 23136 11456
rect 23072 11396 23076 11452
rect 23076 11396 23132 11452
rect 23132 11396 23136 11452
rect 23072 11392 23136 11396
rect 23152 11452 23216 11456
rect 23152 11396 23156 11452
rect 23156 11396 23212 11452
rect 23212 11396 23216 11452
rect 23152 11392 23216 11396
rect 23232 11452 23296 11456
rect 23232 11396 23236 11452
rect 23236 11396 23292 11452
rect 23292 11396 23296 11452
rect 23232 11392 23296 11396
rect 3652 10908 3716 10912
rect 3652 10852 3656 10908
rect 3656 10852 3712 10908
rect 3712 10852 3716 10908
rect 3652 10848 3716 10852
rect 3732 10908 3796 10912
rect 3732 10852 3736 10908
rect 3736 10852 3792 10908
rect 3792 10852 3796 10908
rect 3732 10848 3796 10852
rect 3812 10908 3876 10912
rect 3812 10852 3816 10908
rect 3816 10852 3872 10908
rect 3872 10852 3876 10908
rect 3812 10848 3876 10852
rect 3892 10908 3956 10912
rect 3892 10852 3896 10908
rect 3896 10852 3952 10908
rect 3952 10852 3956 10908
rect 3892 10848 3956 10852
rect 3972 10908 4036 10912
rect 3972 10852 3976 10908
rect 3976 10852 4032 10908
rect 4032 10852 4036 10908
rect 3972 10848 4036 10852
rect 7652 10908 7716 10912
rect 7652 10852 7656 10908
rect 7656 10852 7712 10908
rect 7712 10852 7716 10908
rect 7652 10848 7716 10852
rect 7732 10908 7796 10912
rect 7732 10852 7736 10908
rect 7736 10852 7792 10908
rect 7792 10852 7796 10908
rect 7732 10848 7796 10852
rect 7812 10908 7876 10912
rect 7812 10852 7816 10908
rect 7816 10852 7872 10908
rect 7872 10852 7876 10908
rect 7812 10848 7876 10852
rect 7892 10908 7956 10912
rect 7892 10852 7896 10908
rect 7896 10852 7952 10908
rect 7952 10852 7956 10908
rect 7892 10848 7956 10852
rect 7972 10908 8036 10912
rect 7972 10852 7976 10908
rect 7976 10852 8032 10908
rect 8032 10852 8036 10908
rect 7972 10848 8036 10852
rect 11652 10908 11716 10912
rect 11652 10852 11656 10908
rect 11656 10852 11712 10908
rect 11712 10852 11716 10908
rect 11652 10848 11716 10852
rect 11732 10908 11796 10912
rect 11732 10852 11736 10908
rect 11736 10852 11792 10908
rect 11792 10852 11796 10908
rect 11732 10848 11796 10852
rect 11812 10908 11876 10912
rect 11812 10852 11816 10908
rect 11816 10852 11872 10908
rect 11872 10852 11876 10908
rect 11812 10848 11876 10852
rect 11892 10908 11956 10912
rect 11892 10852 11896 10908
rect 11896 10852 11952 10908
rect 11952 10852 11956 10908
rect 11892 10848 11956 10852
rect 11972 10908 12036 10912
rect 11972 10852 11976 10908
rect 11976 10852 12032 10908
rect 12032 10852 12036 10908
rect 11972 10848 12036 10852
rect 15652 10908 15716 10912
rect 15652 10852 15656 10908
rect 15656 10852 15712 10908
rect 15712 10852 15716 10908
rect 15652 10848 15716 10852
rect 15732 10908 15796 10912
rect 15732 10852 15736 10908
rect 15736 10852 15792 10908
rect 15792 10852 15796 10908
rect 15732 10848 15796 10852
rect 15812 10908 15876 10912
rect 15812 10852 15816 10908
rect 15816 10852 15872 10908
rect 15872 10852 15876 10908
rect 15812 10848 15876 10852
rect 15892 10908 15956 10912
rect 15892 10852 15896 10908
rect 15896 10852 15952 10908
rect 15952 10852 15956 10908
rect 15892 10848 15956 10852
rect 15972 10908 16036 10912
rect 15972 10852 15976 10908
rect 15976 10852 16032 10908
rect 16032 10852 16036 10908
rect 15972 10848 16036 10852
rect 19652 10908 19716 10912
rect 19652 10852 19656 10908
rect 19656 10852 19712 10908
rect 19712 10852 19716 10908
rect 19652 10848 19716 10852
rect 19732 10908 19796 10912
rect 19732 10852 19736 10908
rect 19736 10852 19792 10908
rect 19792 10852 19796 10908
rect 19732 10848 19796 10852
rect 19812 10908 19876 10912
rect 19812 10852 19816 10908
rect 19816 10852 19872 10908
rect 19872 10852 19876 10908
rect 19812 10848 19876 10852
rect 19892 10908 19956 10912
rect 19892 10852 19896 10908
rect 19896 10852 19952 10908
rect 19952 10852 19956 10908
rect 19892 10848 19956 10852
rect 19972 10908 20036 10912
rect 19972 10852 19976 10908
rect 19976 10852 20032 10908
rect 20032 10852 20036 10908
rect 19972 10848 20036 10852
rect 23652 10908 23716 10912
rect 23652 10852 23656 10908
rect 23656 10852 23712 10908
rect 23712 10852 23716 10908
rect 23652 10848 23716 10852
rect 23732 10908 23796 10912
rect 23732 10852 23736 10908
rect 23736 10852 23792 10908
rect 23792 10852 23796 10908
rect 23732 10848 23796 10852
rect 23812 10908 23876 10912
rect 23812 10852 23816 10908
rect 23816 10852 23872 10908
rect 23872 10852 23876 10908
rect 23812 10848 23876 10852
rect 23892 10908 23956 10912
rect 23892 10852 23896 10908
rect 23896 10852 23952 10908
rect 23952 10852 23956 10908
rect 23892 10848 23956 10852
rect 23972 10908 24036 10912
rect 23972 10852 23976 10908
rect 23976 10852 24032 10908
rect 24032 10852 24036 10908
rect 23972 10848 24036 10852
rect 10180 10780 10244 10844
rect 17356 10704 17420 10708
rect 17356 10648 17370 10704
rect 17370 10648 17420 10704
rect 17356 10644 17420 10648
rect 2912 10364 2976 10368
rect 2912 10308 2916 10364
rect 2916 10308 2972 10364
rect 2972 10308 2976 10364
rect 2912 10304 2976 10308
rect 2992 10364 3056 10368
rect 2992 10308 2996 10364
rect 2996 10308 3052 10364
rect 3052 10308 3056 10364
rect 2992 10304 3056 10308
rect 3072 10364 3136 10368
rect 3072 10308 3076 10364
rect 3076 10308 3132 10364
rect 3132 10308 3136 10364
rect 3072 10304 3136 10308
rect 3152 10364 3216 10368
rect 3152 10308 3156 10364
rect 3156 10308 3212 10364
rect 3212 10308 3216 10364
rect 3152 10304 3216 10308
rect 3232 10364 3296 10368
rect 3232 10308 3236 10364
rect 3236 10308 3292 10364
rect 3292 10308 3296 10364
rect 3232 10304 3296 10308
rect 6912 10364 6976 10368
rect 6912 10308 6916 10364
rect 6916 10308 6972 10364
rect 6972 10308 6976 10364
rect 6912 10304 6976 10308
rect 6992 10364 7056 10368
rect 6992 10308 6996 10364
rect 6996 10308 7052 10364
rect 7052 10308 7056 10364
rect 6992 10304 7056 10308
rect 7072 10364 7136 10368
rect 7072 10308 7076 10364
rect 7076 10308 7132 10364
rect 7132 10308 7136 10364
rect 7072 10304 7136 10308
rect 7152 10364 7216 10368
rect 7152 10308 7156 10364
rect 7156 10308 7212 10364
rect 7212 10308 7216 10364
rect 7152 10304 7216 10308
rect 7232 10364 7296 10368
rect 7232 10308 7236 10364
rect 7236 10308 7292 10364
rect 7292 10308 7296 10364
rect 7232 10304 7296 10308
rect 10912 10364 10976 10368
rect 10912 10308 10916 10364
rect 10916 10308 10972 10364
rect 10972 10308 10976 10364
rect 10912 10304 10976 10308
rect 10992 10364 11056 10368
rect 10992 10308 10996 10364
rect 10996 10308 11052 10364
rect 11052 10308 11056 10364
rect 10992 10304 11056 10308
rect 11072 10364 11136 10368
rect 11072 10308 11076 10364
rect 11076 10308 11132 10364
rect 11132 10308 11136 10364
rect 11072 10304 11136 10308
rect 11152 10364 11216 10368
rect 11152 10308 11156 10364
rect 11156 10308 11212 10364
rect 11212 10308 11216 10364
rect 11152 10304 11216 10308
rect 11232 10364 11296 10368
rect 11232 10308 11236 10364
rect 11236 10308 11292 10364
rect 11292 10308 11296 10364
rect 11232 10304 11296 10308
rect 14912 10364 14976 10368
rect 14912 10308 14916 10364
rect 14916 10308 14972 10364
rect 14972 10308 14976 10364
rect 14912 10304 14976 10308
rect 14992 10364 15056 10368
rect 14992 10308 14996 10364
rect 14996 10308 15052 10364
rect 15052 10308 15056 10364
rect 14992 10304 15056 10308
rect 15072 10364 15136 10368
rect 15072 10308 15076 10364
rect 15076 10308 15132 10364
rect 15132 10308 15136 10364
rect 15072 10304 15136 10308
rect 15152 10364 15216 10368
rect 15152 10308 15156 10364
rect 15156 10308 15212 10364
rect 15212 10308 15216 10364
rect 15152 10304 15216 10308
rect 15232 10364 15296 10368
rect 15232 10308 15236 10364
rect 15236 10308 15292 10364
rect 15292 10308 15296 10364
rect 15232 10304 15296 10308
rect 18912 10364 18976 10368
rect 18912 10308 18916 10364
rect 18916 10308 18972 10364
rect 18972 10308 18976 10364
rect 18912 10304 18976 10308
rect 18992 10364 19056 10368
rect 18992 10308 18996 10364
rect 18996 10308 19052 10364
rect 19052 10308 19056 10364
rect 18992 10304 19056 10308
rect 19072 10364 19136 10368
rect 19072 10308 19076 10364
rect 19076 10308 19132 10364
rect 19132 10308 19136 10364
rect 19072 10304 19136 10308
rect 19152 10364 19216 10368
rect 19152 10308 19156 10364
rect 19156 10308 19212 10364
rect 19212 10308 19216 10364
rect 19152 10304 19216 10308
rect 19232 10364 19296 10368
rect 19232 10308 19236 10364
rect 19236 10308 19292 10364
rect 19292 10308 19296 10364
rect 19232 10304 19296 10308
rect 22912 10364 22976 10368
rect 22912 10308 22916 10364
rect 22916 10308 22972 10364
rect 22972 10308 22976 10364
rect 22912 10304 22976 10308
rect 22992 10364 23056 10368
rect 22992 10308 22996 10364
rect 22996 10308 23052 10364
rect 23052 10308 23056 10364
rect 22992 10304 23056 10308
rect 23072 10364 23136 10368
rect 23072 10308 23076 10364
rect 23076 10308 23132 10364
rect 23132 10308 23136 10364
rect 23072 10304 23136 10308
rect 23152 10364 23216 10368
rect 23152 10308 23156 10364
rect 23156 10308 23212 10364
rect 23212 10308 23216 10364
rect 23152 10304 23216 10308
rect 23232 10364 23296 10368
rect 23232 10308 23236 10364
rect 23236 10308 23292 10364
rect 23292 10308 23296 10364
rect 23232 10304 23296 10308
rect 17540 10296 17604 10300
rect 17540 10240 17554 10296
rect 17554 10240 17604 10296
rect 17540 10236 17604 10240
rect 18276 10236 18340 10300
rect 3652 9820 3716 9824
rect 3652 9764 3656 9820
rect 3656 9764 3712 9820
rect 3712 9764 3716 9820
rect 3652 9760 3716 9764
rect 3732 9820 3796 9824
rect 3732 9764 3736 9820
rect 3736 9764 3792 9820
rect 3792 9764 3796 9820
rect 3732 9760 3796 9764
rect 3812 9820 3876 9824
rect 3812 9764 3816 9820
rect 3816 9764 3872 9820
rect 3872 9764 3876 9820
rect 3812 9760 3876 9764
rect 3892 9820 3956 9824
rect 3892 9764 3896 9820
rect 3896 9764 3952 9820
rect 3952 9764 3956 9820
rect 3892 9760 3956 9764
rect 3972 9820 4036 9824
rect 3972 9764 3976 9820
rect 3976 9764 4032 9820
rect 4032 9764 4036 9820
rect 3972 9760 4036 9764
rect 7652 9820 7716 9824
rect 7652 9764 7656 9820
rect 7656 9764 7712 9820
rect 7712 9764 7716 9820
rect 7652 9760 7716 9764
rect 7732 9820 7796 9824
rect 7732 9764 7736 9820
rect 7736 9764 7792 9820
rect 7792 9764 7796 9820
rect 7732 9760 7796 9764
rect 7812 9820 7876 9824
rect 7812 9764 7816 9820
rect 7816 9764 7872 9820
rect 7872 9764 7876 9820
rect 7812 9760 7876 9764
rect 7892 9820 7956 9824
rect 7892 9764 7896 9820
rect 7896 9764 7952 9820
rect 7952 9764 7956 9820
rect 7892 9760 7956 9764
rect 7972 9820 8036 9824
rect 7972 9764 7976 9820
rect 7976 9764 8032 9820
rect 8032 9764 8036 9820
rect 7972 9760 8036 9764
rect 11652 9820 11716 9824
rect 11652 9764 11656 9820
rect 11656 9764 11712 9820
rect 11712 9764 11716 9820
rect 11652 9760 11716 9764
rect 11732 9820 11796 9824
rect 11732 9764 11736 9820
rect 11736 9764 11792 9820
rect 11792 9764 11796 9820
rect 11732 9760 11796 9764
rect 11812 9820 11876 9824
rect 11812 9764 11816 9820
rect 11816 9764 11872 9820
rect 11872 9764 11876 9820
rect 11812 9760 11876 9764
rect 11892 9820 11956 9824
rect 11892 9764 11896 9820
rect 11896 9764 11952 9820
rect 11952 9764 11956 9820
rect 11892 9760 11956 9764
rect 11972 9820 12036 9824
rect 11972 9764 11976 9820
rect 11976 9764 12032 9820
rect 12032 9764 12036 9820
rect 11972 9760 12036 9764
rect 15652 9820 15716 9824
rect 15652 9764 15656 9820
rect 15656 9764 15712 9820
rect 15712 9764 15716 9820
rect 15652 9760 15716 9764
rect 15732 9820 15796 9824
rect 15732 9764 15736 9820
rect 15736 9764 15792 9820
rect 15792 9764 15796 9820
rect 15732 9760 15796 9764
rect 15812 9820 15876 9824
rect 15812 9764 15816 9820
rect 15816 9764 15872 9820
rect 15872 9764 15876 9820
rect 15812 9760 15876 9764
rect 15892 9820 15956 9824
rect 15892 9764 15896 9820
rect 15896 9764 15952 9820
rect 15952 9764 15956 9820
rect 15892 9760 15956 9764
rect 15972 9820 16036 9824
rect 15972 9764 15976 9820
rect 15976 9764 16032 9820
rect 16032 9764 16036 9820
rect 15972 9760 16036 9764
rect 19652 9820 19716 9824
rect 19652 9764 19656 9820
rect 19656 9764 19712 9820
rect 19712 9764 19716 9820
rect 19652 9760 19716 9764
rect 19732 9820 19796 9824
rect 19732 9764 19736 9820
rect 19736 9764 19792 9820
rect 19792 9764 19796 9820
rect 19732 9760 19796 9764
rect 19812 9820 19876 9824
rect 19812 9764 19816 9820
rect 19816 9764 19872 9820
rect 19872 9764 19876 9820
rect 19812 9760 19876 9764
rect 19892 9820 19956 9824
rect 19892 9764 19896 9820
rect 19896 9764 19952 9820
rect 19952 9764 19956 9820
rect 19892 9760 19956 9764
rect 19972 9820 20036 9824
rect 19972 9764 19976 9820
rect 19976 9764 20032 9820
rect 20032 9764 20036 9820
rect 19972 9760 20036 9764
rect 23652 9820 23716 9824
rect 23652 9764 23656 9820
rect 23656 9764 23712 9820
rect 23712 9764 23716 9820
rect 23652 9760 23716 9764
rect 23732 9820 23796 9824
rect 23732 9764 23736 9820
rect 23736 9764 23792 9820
rect 23792 9764 23796 9820
rect 23732 9760 23796 9764
rect 23812 9820 23876 9824
rect 23812 9764 23816 9820
rect 23816 9764 23872 9820
rect 23872 9764 23876 9820
rect 23812 9760 23876 9764
rect 23892 9820 23956 9824
rect 23892 9764 23896 9820
rect 23896 9764 23952 9820
rect 23952 9764 23956 9820
rect 23892 9760 23956 9764
rect 23972 9820 24036 9824
rect 23972 9764 23976 9820
rect 23976 9764 24032 9820
rect 24032 9764 24036 9820
rect 23972 9760 24036 9764
rect 2912 9276 2976 9280
rect 2912 9220 2916 9276
rect 2916 9220 2972 9276
rect 2972 9220 2976 9276
rect 2912 9216 2976 9220
rect 2992 9276 3056 9280
rect 2992 9220 2996 9276
rect 2996 9220 3052 9276
rect 3052 9220 3056 9276
rect 2992 9216 3056 9220
rect 3072 9276 3136 9280
rect 3072 9220 3076 9276
rect 3076 9220 3132 9276
rect 3132 9220 3136 9276
rect 3072 9216 3136 9220
rect 3152 9276 3216 9280
rect 3152 9220 3156 9276
rect 3156 9220 3212 9276
rect 3212 9220 3216 9276
rect 3152 9216 3216 9220
rect 3232 9276 3296 9280
rect 3232 9220 3236 9276
rect 3236 9220 3292 9276
rect 3292 9220 3296 9276
rect 3232 9216 3296 9220
rect 6912 9276 6976 9280
rect 6912 9220 6916 9276
rect 6916 9220 6972 9276
rect 6972 9220 6976 9276
rect 6912 9216 6976 9220
rect 6992 9276 7056 9280
rect 6992 9220 6996 9276
rect 6996 9220 7052 9276
rect 7052 9220 7056 9276
rect 6992 9216 7056 9220
rect 7072 9276 7136 9280
rect 7072 9220 7076 9276
rect 7076 9220 7132 9276
rect 7132 9220 7136 9276
rect 7072 9216 7136 9220
rect 7152 9276 7216 9280
rect 7152 9220 7156 9276
rect 7156 9220 7212 9276
rect 7212 9220 7216 9276
rect 7152 9216 7216 9220
rect 7232 9276 7296 9280
rect 7232 9220 7236 9276
rect 7236 9220 7292 9276
rect 7292 9220 7296 9276
rect 7232 9216 7296 9220
rect 10912 9276 10976 9280
rect 10912 9220 10916 9276
rect 10916 9220 10972 9276
rect 10972 9220 10976 9276
rect 10912 9216 10976 9220
rect 10992 9276 11056 9280
rect 10992 9220 10996 9276
rect 10996 9220 11052 9276
rect 11052 9220 11056 9276
rect 10992 9216 11056 9220
rect 11072 9276 11136 9280
rect 11072 9220 11076 9276
rect 11076 9220 11132 9276
rect 11132 9220 11136 9276
rect 11072 9216 11136 9220
rect 11152 9276 11216 9280
rect 11152 9220 11156 9276
rect 11156 9220 11212 9276
rect 11212 9220 11216 9276
rect 11152 9216 11216 9220
rect 11232 9276 11296 9280
rect 11232 9220 11236 9276
rect 11236 9220 11292 9276
rect 11292 9220 11296 9276
rect 11232 9216 11296 9220
rect 14912 9276 14976 9280
rect 14912 9220 14916 9276
rect 14916 9220 14972 9276
rect 14972 9220 14976 9276
rect 14912 9216 14976 9220
rect 14992 9276 15056 9280
rect 14992 9220 14996 9276
rect 14996 9220 15052 9276
rect 15052 9220 15056 9276
rect 14992 9216 15056 9220
rect 15072 9276 15136 9280
rect 15072 9220 15076 9276
rect 15076 9220 15132 9276
rect 15132 9220 15136 9276
rect 15072 9216 15136 9220
rect 15152 9276 15216 9280
rect 15152 9220 15156 9276
rect 15156 9220 15212 9276
rect 15212 9220 15216 9276
rect 15152 9216 15216 9220
rect 15232 9276 15296 9280
rect 15232 9220 15236 9276
rect 15236 9220 15292 9276
rect 15292 9220 15296 9276
rect 15232 9216 15296 9220
rect 18912 9276 18976 9280
rect 18912 9220 18916 9276
rect 18916 9220 18972 9276
rect 18972 9220 18976 9276
rect 18912 9216 18976 9220
rect 18992 9276 19056 9280
rect 18992 9220 18996 9276
rect 18996 9220 19052 9276
rect 19052 9220 19056 9276
rect 18992 9216 19056 9220
rect 19072 9276 19136 9280
rect 19072 9220 19076 9276
rect 19076 9220 19132 9276
rect 19132 9220 19136 9276
rect 19072 9216 19136 9220
rect 19152 9276 19216 9280
rect 19152 9220 19156 9276
rect 19156 9220 19212 9276
rect 19212 9220 19216 9276
rect 19152 9216 19216 9220
rect 19232 9276 19296 9280
rect 19232 9220 19236 9276
rect 19236 9220 19292 9276
rect 19292 9220 19296 9276
rect 19232 9216 19296 9220
rect 22912 9276 22976 9280
rect 22912 9220 22916 9276
rect 22916 9220 22972 9276
rect 22972 9220 22976 9276
rect 22912 9216 22976 9220
rect 22992 9276 23056 9280
rect 22992 9220 22996 9276
rect 22996 9220 23052 9276
rect 23052 9220 23056 9276
rect 22992 9216 23056 9220
rect 23072 9276 23136 9280
rect 23072 9220 23076 9276
rect 23076 9220 23132 9276
rect 23132 9220 23136 9276
rect 23072 9216 23136 9220
rect 23152 9276 23216 9280
rect 23152 9220 23156 9276
rect 23156 9220 23212 9276
rect 23212 9220 23216 9276
rect 23152 9216 23216 9220
rect 23232 9276 23296 9280
rect 23232 9220 23236 9276
rect 23236 9220 23292 9276
rect 23292 9220 23296 9276
rect 23232 9216 23296 9220
rect 3652 8732 3716 8736
rect 3652 8676 3656 8732
rect 3656 8676 3712 8732
rect 3712 8676 3716 8732
rect 3652 8672 3716 8676
rect 3732 8732 3796 8736
rect 3732 8676 3736 8732
rect 3736 8676 3792 8732
rect 3792 8676 3796 8732
rect 3732 8672 3796 8676
rect 3812 8732 3876 8736
rect 3812 8676 3816 8732
rect 3816 8676 3872 8732
rect 3872 8676 3876 8732
rect 3812 8672 3876 8676
rect 3892 8732 3956 8736
rect 3892 8676 3896 8732
rect 3896 8676 3952 8732
rect 3952 8676 3956 8732
rect 3892 8672 3956 8676
rect 3972 8732 4036 8736
rect 3972 8676 3976 8732
rect 3976 8676 4032 8732
rect 4032 8676 4036 8732
rect 3972 8672 4036 8676
rect 7652 8732 7716 8736
rect 7652 8676 7656 8732
rect 7656 8676 7712 8732
rect 7712 8676 7716 8732
rect 7652 8672 7716 8676
rect 7732 8732 7796 8736
rect 7732 8676 7736 8732
rect 7736 8676 7792 8732
rect 7792 8676 7796 8732
rect 7732 8672 7796 8676
rect 7812 8732 7876 8736
rect 7812 8676 7816 8732
rect 7816 8676 7872 8732
rect 7872 8676 7876 8732
rect 7812 8672 7876 8676
rect 7892 8732 7956 8736
rect 7892 8676 7896 8732
rect 7896 8676 7952 8732
rect 7952 8676 7956 8732
rect 7892 8672 7956 8676
rect 7972 8732 8036 8736
rect 7972 8676 7976 8732
rect 7976 8676 8032 8732
rect 8032 8676 8036 8732
rect 7972 8672 8036 8676
rect 11652 8732 11716 8736
rect 11652 8676 11656 8732
rect 11656 8676 11712 8732
rect 11712 8676 11716 8732
rect 11652 8672 11716 8676
rect 11732 8732 11796 8736
rect 11732 8676 11736 8732
rect 11736 8676 11792 8732
rect 11792 8676 11796 8732
rect 11732 8672 11796 8676
rect 11812 8732 11876 8736
rect 11812 8676 11816 8732
rect 11816 8676 11872 8732
rect 11872 8676 11876 8732
rect 11812 8672 11876 8676
rect 11892 8732 11956 8736
rect 11892 8676 11896 8732
rect 11896 8676 11952 8732
rect 11952 8676 11956 8732
rect 11892 8672 11956 8676
rect 11972 8732 12036 8736
rect 11972 8676 11976 8732
rect 11976 8676 12032 8732
rect 12032 8676 12036 8732
rect 11972 8672 12036 8676
rect 15652 8732 15716 8736
rect 15652 8676 15656 8732
rect 15656 8676 15712 8732
rect 15712 8676 15716 8732
rect 15652 8672 15716 8676
rect 15732 8732 15796 8736
rect 15732 8676 15736 8732
rect 15736 8676 15792 8732
rect 15792 8676 15796 8732
rect 15732 8672 15796 8676
rect 15812 8732 15876 8736
rect 15812 8676 15816 8732
rect 15816 8676 15872 8732
rect 15872 8676 15876 8732
rect 15812 8672 15876 8676
rect 15892 8732 15956 8736
rect 15892 8676 15896 8732
rect 15896 8676 15952 8732
rect 15952 8676 15956 8732
rect 15892 8672 15956 8676
rect 15972 8732 16036 8736
rect 15972 8676 15976 8732
rect 15976 8676 16032 8732
rect 16032 8676 16036 8732
rect 15972 8672 16036 8676
rect 19652 8732 19716 8736
rect 19652 8676 19656 8732
rect 19656 8676 19712 8732
rect 19712 8676 19716 8732
rect 19652 8672 19716 8676
rect 19732 8732 19796 8736
rect 19732 8676 19736 8732
rect 19736 8676 19792 8732
rect 19792 8676 19796 8732
rect 19732 8672 19796 8676
rect 19812 8732 19876 8736
rect 19812 8676 19816 8732
rect 19816 8676 19872 8732
rect 19872 8676 19876 8732
rect 19812 8672 19876 8676
rect 19892 8732 19956 8736
rect 19892 8676 19896 8732
rect 19896 8676 19952 8732
rect 19952 8676 19956 8732
rect 19892 8672 19956 8676
rect 19972 8732 20036 8736
rect 19972 8676 19976 8732
rect 19976 8676 20032 8732
rect 20032 8676 20036 8732
rect 19972 8672 20036 8676
rect 23652 8732 23716 8736
rect 23652 8676 23656 8732
rect 23656 8676 23712 8732
rect 23712 8676 23716 8732
rect 23652 8672 23716 8676
rect 23732 8732 23796 8736
rect 23732 8676 23736 8732
rect 23736 8676 23792 8732
rect 23792 8676 23796 8732
rect 23732 8672 23796 8676
rect 23812 8732 23876 8736
rect 23812 8676 23816 8732
rect 23816 8676 23872 8732
rect 23872 8676 23876 8732
rect 23812 8672 23876 8676
rect 23892 8732 23956 8736
rect 23892 8676 23896 8732
rect 23896 8676 23952 8732
rect 23952 8676 23956 8732
rect 23892 8672 23956 8676
rect 23972 8732 24036 8736
rect 23972 8676 23976 8732
rect 23976 8676 24032 8732
rect 24032 8676 24036 8732
rect 23972 8672 24036 8676
rect 14596 8528 14660 8532
rect 14596 8472 14610 8528
rect 14610 8472 14660 8528
rect 14596 8468 14660 8472
rect 2912 8188 2976 8192
rect 2912 8132 2916 8188
rect 2916 8132 2972 8188
rect 2972 8132 2976 8188
rect 2912 8128 2976 8132
rect 2992 8188 3056 8192
rect 2992 8132 2996 8188
rect 2996 8132 3052 8188
rect 3052 8132 3056 8188
rect 2992 8128 3056 8132
rect 3072 8188 3136 8192
rect 3072 8132 3076 8188
rect 3076 8132 3132 8188
rect 3132 8132 3136 8188
rect 3072 8128 3136 8132
rect 3152 8188 3216 8192
rect 3152 8132 3156 8188
rect 3156 8132 3212 8188
rect 3212 8132 3216 8188
rect 3152 8128 3216 8132
rect 3232 8188 3296 8192
rect 3232 8132 3236 8188
rect 3236 8132 3292 8188
rect 3292 8132 3296 8188
rect 3232 8128 3296 8132
rect 6912 8188 6976 8192
rect 6912 8132 6916 8188
rect 6916 8132 6972 8188
rect 6972 8132 6976 8188
rect 6912 8128 6976 8132
rect 6992 8188 7056 8192
rect 6992 8132 6996 8188
rect 6996 8132 7052 8188
rect 7052 8132 7056 8188
rect 6992 8128 7056 8132
rect 7072 8188 7136 8192
rect 7072 8132 7076 8188
rect 7076 8132 7132 8188
rect 7132 8132 7136 8188
rect 7072 8128 7136 8132
rect 7152 8188 7216 8192
rect 7152 8132 7156 8188
rect 7156 8132 7212 8188
rect 7212 8132 7216 8188
rect 7152 8128 7216 8132
rect 7232 8188 7296 8192
rect 7232 8132 7236 8188
rect 7236 8132 7292 8188
rect 7292 8132 7296 8188
rect 7232 8128 7296 8132
rect 10912 8188 10976 8192
rect 10912 8132 10916 8188
rect 10916 8132 10972 8188
rect 10972 8132 10976 8188
rect 10912 8128 10976 8132
rect 10992 8188 11056 8192
rect 10992 8132 10996 8188
rect 10996 8132 11052 8188
rect 11052 8132 11056 8188
rect 10992 8128 11056 8132
rect 11072 8188 11136 8192
rect 11072 8132 11076 8188
rect 11076 8132 11132 8188
rect 11132 8132 11136 8188
rect 11072 8128 11136 8132
rect 11152 8188 11216 8192
rect 11152 8132 11156 8188
rect 11156 8132 11212 8188
rect 11212 8132 11216 8188
rect 11152 8128 11216 8132
rect 11232 8188 11296 8192
rect 11232 8132 11236 8188
rect 11236 8132 11292 8188
rect 11292 8132 11296 8188
rect 11232 8128 11296 8132
rect 14912 8188 14976 8192
rect 14912 8132 14916 8188
rect 14916 8132 14972 8188
rect 14972 8132 14976 8188
rect 14912 8128 14976 8132
rect 14992 8188 15056 8192
rect 14992 8132 14996 8188
rect 14996 8132 15052 8188
rect 15052 8132 15056 8188
rect 14992 8128 15056 8132
rect 15072 8188 15136 8192
rect 15072 8132 15076 8188
rect 15076 8132 15132 8188
rect 15132 8132 15136 8188
rect 15072 8128 15136 8132
rect 15152 8188 15216 8192
rect 15152 8132 15156 8188
rect 15156 8132 15212 8188
rect 15212 8132 15216 8188
rect 15152 8128 15216 8132
rect 15232 8188 15296 8192
rect 15232 8132 15236 8188
rect 15236 8132 15292 8188
rect 15292 8132 15296 8188
rect 15232 8128 15296 8132
rect 18912 8188 18976 8192
rect 18912 8132 18916 8188
rect 18916 8132 18972 8188
rect 18972 8132 18976 8188
rect 18912 8128 18976 8132
rect 18992 8188 19056 8192
rect 18992 8132 18996 8188
rect 18996 8132 19052 8188
rect 19052 8132 19056 8188
rect 18992 8128 19056 8132
rect 19072 8188 19136 8192
rect 19072 8132 19076 8188
rect 19076 8132 19132 8188
rect 19132 8132 19136 8188
rect 19072 8128 19136 8132
rect 19152 8188 19216 8192
rect 19152 8132 19156 8188
rect 19156 8132 19212 8188
rect 19212 8132 19216 8188
rect 19152 8128 19216 8132
rect 19232 8188 19296 8192
rect 19232 8132 19236 8188
rect 19236 8132 19292 8188
rect 19292 8132 19296 8188
rect 19232 8128 19296 8132
rect 22912 8188 22976 8192
rect 22912 8132 22916 8188
rect 22916 8132 22972 8188
rect 22972 8132 22976 8188
rect 22912 8128 22976 8132
rect 22992 8188 23056 8192
rect 22992 8132 22996 8188
rect 22996 8132 23052 8188
rect 23052 8132 23056 8188
rect 22992 8128 23056 8132
rect 23072 8188 23136 8192
rect 23072 8132 23076 8188
rect 23076 8132 23132 8188
rect 23132 8132 23136 8188
rect 23072 8128 23136 8132
rect 23152 8188 23216 8192
rect 23152 8132 23156 8188
rect 23156 8132 23212 8188
rect 23212 8132 23216 8188
rect 23152 8128 23216 8132
rect 23232 8188 23296 8192
rect 23232 8132 23236 8188
rect 23236 8132 23292 8188
rect 23292 8132 23296 8188
rect 23232 8128 23296 8132
rect 18644 7924 18708 7988
rect 3652 7644 3716 7648
rect 3652 7588 3656 7644
rect 3656 7588 3712 7644
rect 3712 7588 3716 7644
rect 3652 7584 3716 7588
rect 3732 7644 3796 7648
rect 3732 7588 3736 7644
rect 3736 7588 3792 7644
rect 3792 7588 3796 7644
rect 3732 7584 3796 7588
rect 3812 7644 3876 7648
rect 3812 7588 3816 7644
rect 3816 7588 3872 7644
rect 3872 7588 3876 7644
rect 3812 7584 3876 7588
rect 3892 7644 3956 7648
rect 3892 7588 3896 7644
rect 3896 7588 3952 7644
rect 3952 7588 3956 7644
rect 3892 7584 3956 7588
rect 3972 7644 4036 7648
rect 3972 7588 3976 7644
rect 3976 7588 4032 7644
rect 4032 7588 4036 7644
rect 3972 7584 4036 7588
rect 7652 7644 7716 7648
rect 7652 7588 7656 7644
rect 7656 7588 7712 7644
rect 7712 7588 7716 7644
rect 7652 7584 7716 7588
rect 7732 7644 7796 7648
rect 7732 7588 7736 7644
rect 7736 7588 7792 7644
rect 7792 7588 7796 7644
rect 7732 7584 7796 7588
rect 7812 7644 7876 7648
rect 7812 7588 7816 7644
rect 7816 7588 7872 7644
rect 7872 7588 7876 7644
rect 7812 7584 7876 7588
rect 7892 7644 7956 7648
rect 7892 7588 7896 7644
rect 7896 7588 7952 7644
rect 7952 7588 7956 7644
rect 7892 7584 7956 7588
rect 7972 7644 8036 7648
rect 7972 7588 7976 7644
rect 7976 7588 8032 7644
rect 8032 7588 8036 7644
rect 7972 7584 8036 7588
rect 11652 7644 11716 7648
rect 11652 7588 11656 7644
rect 11656 7588 11712 7644
rect 11712 7588 11716 7644
rect 11652 7584 11716 7588
rect 11732 7644 11796 7648
rect 11732 7588 11736 7644
rect 11736 7588 11792 7644
rect 11792 7588 11796 7644
rect 11732 7584 11796 7588
rect 11812 7644 11876 7648
rect 11812 7588 11816 7644
rect 11816 7588 11872 7644
rect 11872 7588 11876 7644
rect 11812 7584 11876 7588
rect 11892 7644 11956 7648
rect 11892 7588 11896 7644
rect 11896 7588 11952 7644
rect 11952 7588 11956 7644
rect 11892 7584 11956 7588
rect 11972 7644 12036 7648
rect 11972 7588 11976 7644
rect 11976 7588 12032 7644
rect 12032 7588 12036 7644
rect 11972 7584 12036 7588
rect 15652 7644 15716 7648
rect 15652 7588 15656 7644
rect 15656 7588 15712 7644
rect 15712 7588 15716 7644
rect 15652 7584 15716 7588
rect 15732 7644 15796 7648
rect 15732 7588 15736 7644
rect 15736 7588 15792 7644
rect 15792 7588 15796 7644
rect 15732 7584 15796 7588
rect 15812 7644 15876 7648
rect 15812 7588 15816 7644
rect 15816 7588 15872 7644
rect 15872 7588 15876 7644
rect 15812 7584 15876 7588
rect 15892 7644 15956 7648
rect 15892 7588 15896 7644
rect 15896 7588 15952 7644
rect 15952 7588 15956 7644
rect 15892 7584 15956 7588
rect 15972 7644 16036 7648
rect 15972 7588 15976 7644
rect 15976 7588 16032 7644
rect 16032 7588 16036 7644
rect 15972 7584 16036 7588
rect 19652 7644 19716 7648
rect 19652 7588 19656 7644
rect 19656 7588 19712 7644
rect 19712 7588 19716 7644
rect 19652 7584 19716 7588
rect 19732 7644 19796 7648
rect 19732 7588 19736 7644
rect 19736 7588 19792 7644
rect 19792 7588 19796 7644
rect 19732 7584 19796 7588
rect 19812 7644 19876 7648
rect 19812 7588 19816 7644
rect 19816 7588 19872 7644
rect 19872 7588 19876 7644
rect 19812 7584 19876 7588
rect 19892 7644 19956 7648
rect 19892 7588 19896 7644
rect 19896 7588 19952 7644
rect 19952 7588 19956 7644
rect 19892 7584 19956 7588
rect 19972 7644 20036 7648
rect 19972 7588 19976 7644
rect 19976 7588 20032 7644
rect 20032 7588 20036 7644
rect 19972 7584 20036 7588
rect 23652 7644 23716 7648
rect 23652 7588 23656 7644
rect 23656 7588 23712 7644
rect 23712 7588 23716 7644
rect 23652 7584 23716 7588
rect 23732 7644 23796 7648
rect 23732 7588 23736 7644
rect 23736 7588 23792 7644
rect 23792 7588 23796 7644
rect 23732 7584 23796 7588
rect 23812 7644 23876 7648
rect 23812 7588 23816 7644
rect 23816 7588 23872 7644
rect 23872 7588 23876 7644
rect 23812 7584 23876 7588
rect 23892 7644 23956 7648
rect 23892 7588 23896 7644
rect 23896 7588 23952 7644
rect 23952 7588 23956 7644
rect 23892 7584 23956 7588
rect 23972 7644 24036 7648
rect 23972 7588 23976 7644
rect 23976 7588 24032 7644
rect 24032 7588 24036 7644
rect 23972 7584 24036 7588
rect 2912 7100 2976 7104
rect 2912 7044 2916 7100
rect 2916 7044 2972 7100
rect 2972 7044 2976 7100
rect 2912 7040 2976 7044
rect 2992 7100 3056 7104
rect 2992 7044 2996 7100
rect 2996 7044 3052 7100
rect 3052 7044 3056 7100
rect 2992 7040 3056 7044
rect 3072 7100 3136 7104
rect 3072 7044 3076 7100
rect 3076 7044 3132 7100
rect 3132 7044 3136 7100
rect 3072 7040 3136 7044
rect 3152 7100 3216 7104
rect 3152 7044 3156 7100
rect 3156 7044 3212 7100
rect 3212 7044 3216 7100
rect 3152 7040 3216 7044
rect 3232 7100 3296 7104
rect 3232 7044 3236 7100
rect 3236 7044 3292 7100
rect 3292 7044 3296 7100
rect 3232 7040 3296 7044
rect 6912 7100 6976 7104
rect 6912 7044 6916 7100
rect 6916 7044 6972 7100
rect 6972 7044 6976 7100
rect 6912 7040 6976 7044
rect 6992 7100 7056 7104
rect 6992 7044 6996 7100
rect 6996 7044 7052 7100
rect 7052 7044 7056 7100
rect 6992 7040 7056 7044
rect 7072 7100 7136 7104
rect 7072 7044 7076 7100
rect 7076 7044 7132 7100
rect 7132 7044 7136 7100
rect 7072 7040 7136 7044
rect 7152 7100 7216 7104
rect 7152 7044 7156 7100
rect 7156 7044 7212 7100
rect 7212 7044 7216 7100
rect 7152 7040 7216 7044
rect 7232 7100 7296 7104
rect 7232 7044 7236 7100
rect 7236 7044 7292 7100
rect 7292 7044 7296 7100
rect 7232 7040 7296 7044
rect 10912 7100 10976 7104
rect 10912 7044 10916 7100
rect 10916 7044 10972 7100
rect 10972 7044 10976 7100
rect 10912 7040 10976 7044
rect 10992 7100 11056 7104
rect 10992 7044 10996 7100
rect 10996 7044 11052 7100
rect 11052 7044 11056 7100
rect 10992 7040 11056 7044
rect 11072 7100 11136 7104
rect 11072 7044 11076 7100
rect 11076 7044 11132 7100
rect 11132 7044 11136 7100
rect 11072 7040 11136 7044
rect 11152 7100 11216 7104
rect 11152 7044 11156 7100
rect 11156 7044 11212 7100
rect 11212 7044 11216 7100
rect 11152 7040 11216 7044
rect 11232 7100 11296 7104
rect 11232 7044 11236 7100
rect 11236 7044 11292 7100
rect 11292 7044 11296 7100
rect 11232 7040 11296 7044
rect 14912 7100 14976 7104
rect 14912 7044 14916 7100
rect 14916 7044 14972 7100
rect 14972 7044 14976 7100
rect 14912 7040 14976 7044
rect 14992 7100 15056 7104
rect 14992 7044 14996 7100
rect 14996 7044 15052 7100
rect 15052 7044 15056 7100
rect 14992 7040 15056 7044
rect 15072 7100 15136 7104
rect 15072 7044 15076 7100
rect 15076 7044 15132 7100
rect 15132 7044 15136 7100
rect 15072 7040 15136 7044
rect 15152 7100 15216 7104
rect 15152 7044 15156 7100
rect 15156 7044 15212 7100
rect 15212 7044 15216 7100
rect 15152 7040 15216 7044
rect 15232 7100 15296 7104
rect 15232 7044 15236 7100
rect 15236 7044 15292 7100
rect 15292 7044 15296 7100
rect 15232 7040 15296 7044
rect 18912 7100 18976 7104
rect 18912 7044 18916 7100
rect 18916 7044 18972 7100
rect 18972 7044 18976 7100
rect 18912 7040 18976 7044
rect 18992 7100 19056 7104
rect 18992 7044 18996 7100
rect 18996 7044 19052 7100
rect 19052 7044 19056 7100
rect 18992 7040 19056 7044
rect 19072 7100 19136 7104
rect 19072 7044 19076 7100
rect 19076 7044 19132 7100
rect 19132 7044 19136 7100
rect 19072 7040 19136 7044
rect 19152 7100 19216 7104
rect 19152 7044 19156 7100
rect 19156 7044 19212 7100
rect 19212 7044 19216 7100
rect 19152 7040 19216 7044
rect 19232 7100 19296 7104
rect 19232 7044 19236 7100
rect 19236 7044 19292 7100
rect 19292 7044 19296 7100
rect 19232 7040 19296 7044
rect 22912 7100 22976 7104
rect 22912 7044 22916 7100
rect 22916 7044 22972 7100
rect 22972 7044 22976 7100
rect 22912 7040 22976 7044
rect 22992 7100 23056 7104
rect 22992 7044 22996 7100
rect 22996 7044 23052 7100
rect 23052 7044 23056 7100
rect 22992 7040 23056 7044
rect 23072 7100 23136 7104
rect 23072 7044 23076 7100
rect 23076 7044 23132 7100
rect 23132 7044 23136 7100
rect 23072 7040 23136 7044
rect 23152 7100 23216 7104
rect 23152 7044 23156 7100
rect 23156 7044 23212 7100
rect 23212 7044 23216 7100
rect 23152 7040 23216 7044
rect 23232 7100 23296 7104
rect 23232 7044 23236 7100
rect 23236 7044 23292 7100
rect 23292 7044 23296 7100
rect 23232 7040 23296 7044
rect 5212 7032 5276 7036
rect 5212 6976 5226 7032
rect 5226 6976 5276 7032
rect 5212 6972 5276 6976
rect 18460 6700 18524 6764
rect 3652 6556 3716 6560
rect 3652 6500 3656 6556
rect 3656 6500 3712 6556
rect 3712 6500 3716 6556
rect 3652 6496 3716 6500
rect 3732 6556 3796 6560
rect 3732 6500 3736 6556
rect 3736 6500 3792 6556
rect 3792 6500 3796 6556
rect 3732 6496 3796 6500
rect 3812 6556 3876 6560
rect 3812 6500 3816 6556
rect 3816 6500 3872 6556
rect 3872 6500 3876 6556
rect 3812 6496 3876 6500
rect 3892 6556 3956 6560
rect 3892 6500 3896 6556
rect 3896 6500 3952 6556
rect 3952 6500 3956 6556
rect 3892 6496 3956 6500
rect 3972 6556 4036 6560
rect 3972 6500 3976 6556
rect 3976 6500 4032 6556
rect 4032 6500 4036 6556
rect 3972 6496 4036 6500
rect 7652 6556 7716 6560
rect 7652 6500 7656 6556
rect 7656 6500 7712 6556
rect 7712 6500 7716 6556
rect 7652 6496 7716 6500
rect 7732 6556 7796 6560
rect 7732 6500 7736 6556
rect 7736 6500 7792 6556
rect 7792 6500 7796 6556
rect 7732 6496 7796 6500
rect 7812 6556 7876 6560
rect 7812 6500 7816 6556
rect 7816 6500 7872 6556
rect 7872 6500 7876 6556
rect 7812 6496 7876 6500
rect 7892 6556 7956 6560
rect 7892 6500 7896 6556
rect 7896 6500 7952 6556
rect 7952 6500 7956 6556
rect 7892 6496 7956 6500
rect 7972 6556 8036 6560
rect 7972 6500 7976 6556
rect 7976 6500 8032 6556
rect 8032 6500 8036 6556
rect 7972 6496 8036 6500
rect 11652 6556 11716 6560
rect 11652 6500 11656 6556
rect 11656 6500 11712 6556
rect 11712 6500 11716 6556
rect 11652 6496 11716 6500
rect 11732 6556 11796 6560
rect 11732 6500 11736 6556
rect 11736 6500 11792 6556
rect 11792 6500 11796 6556
rect 11732 6496 11796 6500
rect 11812 6556 11876 6560
rect 11812 6500 11816 6556
rect 11816 6500 11872 6556
rect 11872 6500 11876 6556
rect 11812 6496 11876 6500
rect 11892 6556 11956 6560
rect 11892 6500 11896 6556
rect 11896 6500 11952 6556
rect 11952 6500 11956 6556
rect 11892 6496 11956 6500
rect 11972 6556 12036 6560
rect 11972 6500 11976 6556
rect 11976 6500 12032 6556
rect 12032 6500 12036 6556
rect 11972 6496 12036 6500
rect 15652 6556 15716 6560
rect 15652 6500 15656 6556
rect 15656 6500 15712 6556
rect 15712 6500 15716 6556
rect 15652 6496 15716 6500
rect 15732 6556 15796 6560
rect 15732 6500 15736 6556
rect 15736 6500 15792 6556
rect 15792 6500 15796 6556
rect 15732 6496 15796 6500
rect 15812 6556 15876 6560
rect 15812 6500 15816 6556
rect 15816 6500 15872 6556
rect 15872 6500 15876 6556
rect 15812 6496 15876 6500
rect 15892 6556 15956 6560
rect 15892 6500 15896 6556
rect 15896 6500 15952 6556
rect 15952 6500 15956 6556
rect 15892 6496 15956 6500
rect 15972 6556 16036 6560
rect 15972 6500 15976 6556
rect 15976 6500 16032 6556
rect 16032 6500 16036 6556
rect 15972 6496 16036 6500
rect 19652 6556 19716 6560
rect 19652 6500 19656 6556
rect 19656 6500 19712 6556
rect 19712 6500 19716 6556
rect 19652 6496 19716 6500
rect 19732 6556 19796 6560
rect 19732 6500 19736 6556
rect 19736 6500 19792 6556
rect 19792 6500 19796 6556
rect 19732 6496 19796 6500
rect 19812 6556 19876 6560
rect 19812 6500 19816 6556
rect 19816 6500 19872 6556
rect 19872 6500 19876 6556
rect 19812 6496 19876 6500
rect 19892 6556 19956 6560
rect 19892 6500 19896 6556
rect 19896 6500 19952 6556
rect 19952 6500 19956 6556
rect 19892 6496 19956 6500
rect 19972 6556 20036 6560
rect 19972 6500 19976 6556
rect 19976 6500 20032 6556
rect 20032 6500 20036 6556
rect 19972 6496 20036 6500
rect 23652 6556 23716 6560
rect 23652 6500 23656 6556
rect 23656 6500 23712 6556
rect 23712 6500 23716 6556
rect 23652 6496 23716 6500
rect 23732 6556 23796 6560
rect 23732 6500 23736 6556
rect 23736 6500 23792 6556
rect 23792 6500 23796 6556
rect 23732 6496 23796 6500
rect 23812 6556 23876 6560
rect 23812 6500 23816 6556
rect 23816 6500 23872 6556
rect 23872 6500 23876 6556
rect 23812 6496 23876 6500
rect 23892 6556 23956 6560
rect 23892 6500 23896 6556
rect 23896 6500 23952 6556
rect 23952 6500 23956 6556
rect 23892 6496 23956 6500
rect 23972 6556 24036 6560
rect 23972 6500 23976 6556
rect 23976 6500 24032 6556
rect 24032 6500 24036 6556
rect 23972 6496 24036 6500
rect 2912 6012 2976 6016
rect 2912 5956 2916 6012
rect 2916 5956 2972 6012
rect 2972 5956 2976 6012
rect 2912 5952 2976 5956
rect 2992 6012 3056 6016
rect 2992 5956 2996 6012
rect 2996 5956 3052 6012
rect 3052 5956 3056 6012
rect 2992 5952 3056 5956
rect 3072 6012 3136 6016
rect 3072 5956 3076 6012
rect 3076 5956 3132 6012
rect 3132 5956 3136 6012
rect 3072 5952 3136 5956
rect 3152 6012 3216 6016
rect 3152 5956 3156 6012
rect 3156 5956 3212 6012
rect 3212 5956 3216 6012
rect 3152 5952 3216 5956
rect 3232 6012 3296 6016
rect 3232 5956 3236 6012
rect 3236 5956 3292 6012
rect 3292 5956 3296 6012
rect 3232 5952 3296 5956
rect 6912 6012 6976 6016
rect 6912 5956 6916 6012
rect 6916 5956 6972 6012
rect 6972 5956 6976 6012
rect 6912 5952 6976 5956
rect 6992 6012 7056 6016
rect 6992 5956 6996 6012
rect 6996 5956 7052 6012
rect 7052 5956 7056 6012
rect 6992 5952 7056 5956
rect 7072 6012 7136 6016
rect 7072 5956 7076 6012
rect 7076 5956 7132 6012
rect 7132 5956 7136 6012
rect 7072 5952 7136 5956
rect 7152 6012 7216 6016
rect 7152 5956 7156 6012
rect 7156 5956 7212 6012
rect 7212 5956 7216 6012
rect 7152 5952 7216 5956
rect 7232 6012 7296 6016
rect 7232 5956 7236 6012
rect 7236 5956 7292 6012
rect 7292 5956 7296 6012
rect 7232 5952 7296 5956
rect 10912 6012 10976 6016
rect 10912 5956 10916 6012
rect 10916 5956 10972 6012
rect 10972 5956 10976 6012
rect 10912 5952 10976 5956
rect 10992 6012 11056 6016
rect 10992 5956 10996 6012
rect 10996 5956 11052 6012
rect 11052 5956 11056 6012
rect 10992 5952 11056 5956
rect 11072 6012 11136 6016
rect 11072 5956 11076 6012
rect 11076 5956 11132 6012
rect 11132 5956 11136 6012
rect 11072 5952 11136 5956
rect 11152 6012 11216 6016
rect 11152 5956 11156 6012
rect 11156 5956 11212 6012
rect 11212 5956 11216 6012
rect 11152 5952 11216 5956
rect 11232 6012 11296 6016
rect 11232 5956 11236 6012
rect 11236 5956 11292 6012
rect 11292 5956 11296 6012
rect 11232 5952 11296 5956
rect 14912 6012 14976 6016
rect 14912 5956 14916 6012
rect 14916 5956 14972 6012
rect 14972 5956 14976 6012
rect 14912 5952 14976 5956
rect 14992 6012 15056 6016
rect 14992 5956 14996 6012
rect 14996 5956 15052 6012
rect 15052 5956 15056 6012
rect 14992 5952 15056 5956
rect 15072 6012 15136 6016
rect 15072 5956 15076 6012
rect 15076 5956 15132 6012
rect 15132 5956 15136 6012
rect 15072 5952 15136 5956
rect 15152 6012 15216 6016
rect 15152 5956 15156 6012
rect 15156 5956 15212 6012
rect 15212 5956 15216 6012
rect 15152 5952 15216 5956
rect 15232 6012 15296 6016
rect 15232 5956 15236 6012
rect 15236 5956 15292 6012
rect 15292 5956 15296 6012
rect 15232 5952 15296 5956
rect 18912 6012 18976 6016
rect 18912 5956 18916 6012
rect 18916 5956 18972 6012
rect 18972 5956 18976 6012
rect 18912 5952 18976 5956
rect 18992 6012 19056 6016
rect 18992 5956 18996 6012
rect 18996 5956 19052 6012
rect 19052 5956 19056 6012
rect 18992 5952 19056 5956
rect 19072 6012 19136 6016
rect 19072 5956 19076 6012
rect 19076 5956 19132 6012
rect 19132 5956 19136 6012
rect 19072 5952 19136 5956
rect 19152 6012 19216 6016
rect 19152 5956 19156 6012
rect 19156 5956 19212 6012
rect 19212 5956 19216 6012
rect 19152 5952 19216 5956
rect 19232 6012 19296 6016
rect 19232 5956 19236 6012
rect 19236 5956 19292 6012
rect 19292 5956 19296 6012
rect 19232 5952 19296 5956
rect 22912 6012 22976 6016
rect 22912 5956 22916 6012
rect 22916 5956 22972 6012
rect 22972 5956 22976 6012
rect 22912 5952 22976 5956
rect 22992 6012 23056 6016
rect 22992 5956 22996 6012
rect 22996 5956 23052 6012
rect 23052 5956 23056 6012
rect 22992 5952 23056 5956
rect 23072 6012 23136 6016
rect 23072 5956 23076 6012
rect 23076 5956 23132 6012
rect 23132 5956 23136 6012
rect 23072 5952 23136 5956
rect 23152 6012 23216 6016
rect 23152 5956 23156 6012
rect 23156 5956 23212 6012
rect 23212 5956 23216 6012
rect 23152 5952 23216 5956
rect 23232 6012 23296 6016
rect 23232 5956 23236 6012
rect 23236 5956 23292 6012
rect 23292 5956 23296 6012
rect 23232 5952 23296 5956
rect 3652 5468 3716 5472
rect 3652 5412 3656 5468
rect 3656 5412 3712 5468
rect 3712 5412 3716 5468
rect 3652 5408 3716 5412
rect 3732 5468 3796 5472
rect 3732 5412 3736 5468
rect 3736 5412 3792 5468
rect 3792 5412 3796 5468
rect 3732 5408 3796 5412
rect 3812 5468 3876 5472
rect 3812 5412 3816 5468
rect 3816 5412 3872 5468
rect 3872 5412 3876 5468
rect 3812 5408 3876 5412
rect 3892 5468 3956 5472
rect 3892 5412 3896 5468
rect 3896 5412 3952 5468
rect 3952 5412 3956 5468
rect 3892 5408 3956 5412
rect 3972 5468 4036 5472
rect 3972 5412 3976 5468
rect 3976 5412 4032 5468
rect 4032 5412 4036 5468
rect 3972 5408 4036 5412
rect 7652 5468 7716 5472
rect 7652 5412 7656 5468
rect 7656 5412 7712 5468
rect 7712 5412 7716 5468
rect 7652 5408 7716 5412
rect 7732 5468 7796 5472
rect 7732 5412 7736 5468
rect 7736 5412 7792 5468
rect 7792 5412 7796 5468
rect 7732 5408 7796 5412
rect 7812 5468 7876 5472
rect 7812 5412 7816 5468
rect 7816 5412 7872 5468
rect 7872 5412 7876 5468
rect 7812 5408 7876 5412
rect 7892 5468 7956 5472
rect 7892 5412 7896 5468
rect 7896 5412 7952 5468
rect 7952 5412 7956 5468
rect 7892 5408 7956 5412
rect 7972 5468 8036 5472
rect 7972 5412 7976 5468
rect 7976 5412 8032 5468
rect 8032 5412 8036 5468
rect 7972 5408 8036 5412
rect 11652 5468 11716 5472
rect 11652 5412 11656 5468
rect 11656 5412 11712 5468
rect 11712 5412 11716 5468
rect 11652 5408 11716 5412
rect 11732 5468 11796 5472
rect 11732 5412 11736 5468
rect 11736 5412 11792 5468
rect 11792 5412 11796 5468
rect 11732 5408 11796 5412
rect 11812 5468 11876 5472
rect 11812 5412 11816 5468
rect 11816 5412 11872 5468
rect 11872 5412 11876 5468
rect 11812 5408 11876 5412
rect 11892 5468 11956 5472
rect 11892 5412 11896 5468
rect 11896 5412 11952 5468
rect 11952 5412 11956 5468
rect 11892 5408 11956 5412
rect 11972 5468 12036 5472
rect 11972 5412 11976 5468
rect 11976 5412 12032 5468
rect 12032 5412 12036 5468
rect 11972 5408 12036 5412
rect 15652 5468 15716 5472
rect 15652 5412 15656 5468
rect 15656 5412 15712 5468
rect 15712 5412 15716 5468
rect 15652 5408 15716 5412
rect 15732 5468 15796 5472
rect 15732 5412 15736 5468
rect 15736 5412 15792 5468
rect 15792 5412 15796 5468
rect 15732 5408 15796 5412
rect 15812 5468 15876 5472
rect 15812 5412 15816 5468
rect 15816 5412 15872 5468
rect 15872 5412 15876 5468
rect 15812 5408 15876 5412
rect 15892 5468 15956 5472
rect 15892 5412 15896 5468
rect 15896 5412 15952 5468
rect 15952 5412 15956 5468
rect 15892 5408 15956 5412
rect 15972 5468 16036 5472
rect 15972 5412 15976 5468
rect 15976 5412 16032 5468
rect 16032 5412 16036 5468
rect 15972 5408 16036 5412
rect 19652 5468 19716 5472
rect 19652 5412 19656 5468
rect 19656 5412 19712 5468
rect 19712 5412 19716 5468
rect 19652 5408 19716 5412
rect 19732 5468 19796 5472
rect 19732 5412 19736 5468
rect 19736 5412 19792 5468
rect 19792 5412 19796 5468
rect 19732 5408 19796 5412
rect 19812 5468 19876 5472
rect 19812 5412 19816 5468
rect 19816 5412 19872 5468
rect 19872 5412 19876 5468
rect 19812 5408 19876 5412
rect 19892 5468 19956 5472
rect 19892 5412 19896 5468
rect 19896 5412 19952 5468
rect 19952 5412 19956 5468
rect 19892 5408 19956 5412
rect 19972 5468 20036 5472
rect 19972 5412 19976 5468
rect 19976 5412 20032 5468
rect 20032 5412 20036 5468
rect 19972 5408 20036 5412
rect 23652 5468 23716 5472
rect 23652 5412 23656 5468
rect 23656 5412 23712 5468
rect 23712 5412 23716 5468
rect 23652 5408 23716 5412
rect 23732 5468 23796 5472
rect 23732 5412 23736 5468
rect 23736 5412 23792 5468
rect 23792 5412 23796 5468
rect 23732 5408 23796 5412
rect 23812 5468 23876 5472
rect 23812 5412 23816 5468
rect 23816 5412 23872 5468
rect 23872 5412 23876 5468
rect 23812 5408 23876 5412
rect 23892 5468 23956 5472
rect 23892 5412 23896 5468
rect 23896 5412 23952 5468
rect 23952 5412 23956 5468
rect 23892 5408 23956 5412
rect 23972 5468 24036 5472
rect 23972 5412 23976 5468
rect 23976 5412 24032 5468
rect 24032 5412 24036 5468
rect 23972 5408 24036 5412
rect 2912 4924 2976 4928
rect 2912 4868 2916 4924
rect 2916 4868 2972 4924
rect 2972 4868 2976 4924
rect 2912 4864 2976 4868
rect 2992 4924 3056 4928
rect 2992 4868 2996 4924
rect 2996 4868 3052 4924
rect 3052 4868 3056 4924
rect 2992 4864 3056 4868
rect 3072 4924 3136 4928
rect 3072 4868 3076 4924
rect 3076 4868 3132 4924
rect 3132 4868 3136 4924
rect 3072 4864 3136 4868
rect 3152 4924 3216 4928
rect 3152 4868 3156 4924
rect 3156 4868 3212 4924
rect 3212 4868 3216 4924
rect 3152 4864 3216 4868
rect 3232 4924 3296 4928
rect 3232 4868 3236 4924
rect 3236 4868 3292 4924
rect 3292 4868 3296 4924
rect 3232 4864 3296 4868
rect 6912 4924 6976 4928
rect 6912 4868 6916 4924
rect 6916 4868 6972 4924
rect 6972 4868 6976 4924
rect 6912 4864 6976 4868
rect 6992 4924 7056 4928
rect 6992 4868 6996 4924
rect 6996 4868 7052 4924
rect 7052 4868 7056 4924
rect 6992 4864 7056 4868
rect 7072 4924 7136 4928
rect 7072 4868 7076 4924
rect 7076 4868 7132 4924
rect 7132 4868 7136 4924
rect 7072 4864 7136 4868
rect 7152 4924 7216 4928
rect 7152 4868 7156 4924
rect 7156 4868 7212 4924
rect 7212 4868 7216 4924
rect 7152 4864 7216 4868
rect 7232 4924 7296 4928
rect 7232 4868 7236 4924
rect 7236 4868 7292 4924
rect 7292 4868 7296 4924
rect 7232 4864 7296 4868
rect 10912 4924 10976 4928
rect 10912 4868 10916 4924
rect 10916 4868 10972 4924
rect 10972 4868 10976 4924
rect 10912 4864 10976 4868
rect 10992 4924 11056 4928
rect 10992 4868 10996 4924
rect 10996 4868 11052 4924
rect 11052 4868 11056 4924
rect 10992 4864 11056 4868
rect 11072 4924 11136 4928
rect 11072 4868 11076 4924
rect 11076 4868 11132 4924
rect 11132 4868 11136 4924
rect 11072 4864 11136 4868
rect 11152 4924 11216 4928
rect 11152 4868 11156 4924
rect 11156 4868 11212 4924
rect 11212 4868 11216 4924
rect 11152 4864 11216 4868
rect 11232 4924 11296 4928
rect 11232 4868 11236 4924
rect 11236 4868 11292 4924
rect 11292 4868 11296 4924
rect 11232 4864 11296 4868
rect 14912 4924 14976 4928
rect 14912 4868 14916 4924
rect 14916 4868 14972 4924
rect 14972 4868 14976 4924
rect 14912 4864 14976 4868
rect 14992 4924 15056 4928
rect 14992 4868 14996 4924
rect 14996 4868 15052 4924
rect 15052 4868 15056 4924
rect 14992 4864 15056 4868
rect 15072 4924 15136 4928
rect 15072 4868 15076 4924
rect 15076 4868 15132 4924
rect 15132 4868 15136 4924
rect 15072 4864 15136 4868
rect 15152 4924 15216 4928
rect 15152 4868 15156 4924
rect 15156 4868 15212 4924
rect 15212 4868 15216 4924
rect 15152 4864 15216 4868
rect 15232 4924 15296 4928
rect 15232 4868 15236 4924
rect 15236 4868 15292 4924
rect 15292 4868 15296 4924
rect 15232 4864 15296 4868
rect 18912 4924 18976 4928
rect 18912 4868 18916 4924
rect 18916 4868 18972 4924
rect 18972 4868 18976 4924
rect 18912 4864 18976 4868
rect 18992 4924 19056 4928
rect 18992 4868 18996 4924
rect 18996 4868 19052 4924
rect 19052 4868 19056 4924
rect 18992 4864 19056 4868
rect 19072 4924 19136 4928
rect 19072 4868 19076 4924
rect 19076 4868 19132 4924
rect 19132 4868 19136 4924
rect 19072 4864 19136 4868
rect 19152 4924 19216 4928
rect 19152 4868 19156 4924
rect 19156 4868 19212 4924
rect 19212 4868 19216 4924
rect 19152 4864 19216 4868
rect 19232 4924 19296 4928
rect 19232 4868 19236 4924
rect 19236 4868 19292 4924
rect 19292 4868 19296 4924
rect 19232 4864 19296 4868
rect 22912 4924 22976 4928
rect 22912 4868 22916 4924
rect 22916 4868 22972 4924
rect 22972 4868 22976 4924
rect 22912 4864 22976 4868
rect 22992 4924 23056 4928
rect 22992 4868 22996 4924
rect 22996 4868 23052 4924
rect 23052 4868 23056 4924
rect 22992 4864 23056 4868
rect 23072 4924 23136 4928
rect 23072 4868 23076 4924
rect 23076 4868 23132 4924
rect 23132 4868 23136 4924
rect 23072 4864 23136 4868
rect 23152 4924 23216 4928
rect 23152 4868 23156 4924
rect 23156 4868 23212 4924
rect 23212 4868 23216 4924
rect 23152 4864 23216 4868
rect 23232 4924 23296 4928
rect 23232 4868 23236 4924
rect 23236 4868 23292 4924
rect 23292 4868 23296 4924
rect 23232 4864 23296 4868
rect 3652 4380 3716 4384
rect 3652 4324 3656 4380
rect 3656 4324 3712 4380
rect 3712 4324 3716 4380
rect 3652 4320 3716 4324
rect 3732 4380 3796 4384
rect 3732 4324 3736 4380
rect 3736 4324 3792 4380
rect 3792 4324 3796 4380
rect 3732 4320 3796 4324
rect 3812 4380 3876 4384
rect 3812 4324 3816 4380
rect 3816 4324 3872 4380
rect 3872 4324 3876 4380
rect 3812 4320 3876 4324
rect 3892 4380 3956 4384
rect 3892 4324 3896 4380
rect 3896 4324 3952 4380
rect 3952 4324 3956 4380
rect 3892 4320 3956 4324
rect 3972 4380 4036 4384
rect 3972 4324 3976 4380
rect 3976 4324 4032 4380
rect 4032 4324 4036 4380
rect 3972 4320 4036 4324
rect 7652 4380 7716 4384
rect 7652 4324 7656 4380
rect 7656 4324 7712 4380
rect 7712 4324 7716 4380
rect 7652 4320 7716 4324
rect 7732 4380 7796 4384
rect 7732 4324 7736 4380
rect 7736 4324 7792 4380
rect 7792 4324 7796 4380
rect 7732 4320 7796 4324
rect 7812 4380 7876 4384
rect 7812 4324 7816 4380
rect 7816 4324 7872 4380
rect 7872 4324 7876 4380
rect 7812 4320 7876 4324
rect 7892 4380 7956 4384
rect 7892 4324 7896 4380
rect 7896 4324 7952 4380
rect 7952 4324 7956 4380
rect 7892 4320 7956 4324
rect 7972 4380 8036 4384
rect 7972 4324 7976 4380
rect 7976 4324 8032 4380
rect 8032 4324 8036 4380
rect 7972 4320 8036 4324
rect 11652 4380 11716 4384
rect 11652 4324 11656 4380
rect 11656 4324 11712 4380
rect 11712 4324 11716 4380
rect 11652 4320 11716 4324
rect 11732 4380 11796 4384
rect 11732 4324 11736 4380
rect 11736 4324 11792 4380
rect 11792 4324 11796 4380
rect 11732 4320 11796 4324
rect 11812 4380 11876 4384
rect 11812 4324 11816 4380
rect 11816 4324 11872 4380
rect 11872 4324 11876 4380
rect 11812 4320 11876 4324
rect 11892 4380 11956 4384
rect 11892 4324 11896 4380
rect 11896 4324 11952 4380
rect 11952 4324 11956 4380
rect 11892 4320 11956 4324
rect 11972 4380 12036 4384
rect 11972 4324 11976 4380
rect 11976 4324 12032 4380
rect 12032 4324 12036 4380
rect 11972 4320 12036 4324
rect 15652 4380 15716 4384
rect 15652 4324 15656 4380
rect 15656 4324 15712 4380
rect 15712 4324 15716 4380
rect 15652 4320 15716 4324
rect 15732 4380 15796 4384
rect 15732 4324 15736 4380
rect 15736 4324 15792 4380
rect 15792 4324 15796 4380
rect 15732 4320 15796 4324
rect 15812 4380 15876 4384
rect 15812 4324 15816 4380
rect 15816 4324 15872 4380
rect 15872 4324 15876 4380
rect 15812 4320 15876 4324
rect 15892 4380 15956 4384
rect 15892 4324 15896 4380
rect 15896 4324 15952 4380
rect 15952 4324 15956 4380
rect 15892 4320 15956 4324
rect 15972 4380 16036 4384
rect 15972 4324 15976 4380
rect 15976 4324 16032 4380
rect 16032 4324 16036 4380
rect 15972 4320 16036 4324
rect 19652 4380 19716 4384
rect 19652 4324 19656 4380
rect 19656 4324 19712 4380
rect 19712 4324 19716 4380
rect 19652 4320 19716 4324
rect 19732 4380 19796 4384
rect 19732 4324 19736 4380
rect 19736 4324 19792 4380
rect 19792 4324 19796 4380
rect 19732 4320 19796 4324
rect 19812 4380 19876 4384
rect 19812 4324 19816 4380
rect 19816 4324 19872 4380
rect 19872 4324 19876 4380
rect 19812 4320 19876 4324
rect 19892 4380 19956 4384
rect 19892 4324 19896 4380
rect 19896 4324 19952 4380
rect 19952 4324 19956 4380
rect 19892 4320 19956 4324
rect 19972 4380 20036 4384
rect 19972 4324 19976 4380
rect 19976 4324 20032 4380
rect 20032 4324 20036 4380
rect 19972 4320 20036 4324
rect 23652 4380 23716 4384
rect 23652 4324 23656 4380
rect 23656 4324 23712 4380
rect 23712 4324 23716 4380
rect 23652 4320 23716 4324
rect 23732 4380 23796 4384
rect 23732 4324 23736 4380
rect 23736 4324 23792 4380
rect 23792 4324 23796 4380
rect 23732 4320 23796 4324
rect 23812 4380 23876 4384
rect 23812 4324 23816 4380
rect 23816 4324 23872 4380
rect 23872 4324 23876 4380
rect 23812 4320 23876 4324
rect 23892 4380 23956 4384
rect 23892 4324 23896 4380
rect 23896 4324 23952 4380
rect 23952 4324 23956 4380
rect 23892 4320 23956 4324
rect 23972 4380 24036 4384
rect 23972 4324 23976 4380
rect 23976 4324 24032 4380
rect 24032 4324 24036 4380
rect 23972 4320 24036 4324
rect 2912 3836 2976 3840
rect 2912 3780 2916 3836
rect 2916 3780 2972 3836
rect 2972 3780 2976 3836
rect 2912 3776 2976 3780
rect 2992 3836 3056 3840
rect 2992 3780 2996 3836
rect 2996 3780 3052 3836
rect 3052 3780 3056 3836
rect 2992 3776 3056 3780
rect 3072 3836 3136 3840
rect 3072 3780 3076 3836
rect 3076 3780 3132 3836
rect 3132 3780 3136 3836
rect 3072 3776 3136 3780
rect 3152 3836 3216 3840
rect 3152 3780 3156 3836
rect 3156 3780 3212 3836
rect 3212 3780 3216 3836
rect 3152 3776 3216 3780
rect 3232 3836 3296 3840
rect 3232 3780 3236 3836
rect 3236 3780 3292 3836
rect 3292 3780 3296 3836
rect 3232 3776 3296 3780
rect 6912 3836 6976 3840
rect 6912 3780 6916 3836
rect 6916 3780 6972 3836
rect 6972 3780 6976 3836
rect 6912 3776 6976 3780
rect 6992 3836 7056 3840
rect 6992 3780 6996 3836
rect 6996 3780 7052 3836
rect 7052 3780 7056 3836
rect 6992 3776 7056 3780
rect 7072 3836 7136 3840
rect 7072 3780 7076 3836
rect 7076 3780 7132 3836
rect 7132 3780 7136 3836
rect 7072 3776 7136 3780
rect 7152 3836 7216 3840
rect 7152 3780 7156 3836
rect 7156 3780 7212 3836
rect 7212 3780 7216 3836
rect 7152 3776 7216 3780
rect 7232 3836 7296 3840
rect 7232 3780 7236 3836
rect 7236 3780 7292 3836
rect 7292 3780 7296 3836
rect 7232 3776 7296 3780
rect 10912 3836 10976 3840
rect 10912 3780 10916 3836
rect 10916 3780 10972 3836
rect 10972 3780 10976 3836
rect 10912 3776 10976 3780
rect 10992 3836 11056 3840
rect 10992 3780 10996 3836
rect 10996 3780 11052 3836
rect 11052 3780 11056 3836
rect 10992 3776 11056 3780
rect 11072 3836 11136 3840
rect 11072 3780 11076 3836
rect 11076 3780 11132 3836
rect 11132 3780 11136 3836
rect 11072 3776 11136 3780
rect 11152 3836 11216 3840
rect 11152 3780 11156 3836
rect 11156 3780 11212 3836
rect 11212 3780 11216 3836
rect 11152 3776 11216 3780
rect 11232 3836 11296 3840
rect 11232 3780 11236 3836
rect 11236 3780 11292 3836
rect 11292 3780 11296 3836
rect 11232 3776 11296 3780
rect 14912 3836 14976 3840
rect 14912 3780 14916 3836
rect 14916 3780 14972 3836
rect 14972 3780 14976 3836
rect 14912 3776 14976 3780
rect 14992 3836 15056 3840
rect 14992 3780 14996 3836
rect 14996 3780 15052 3836
rect 15052 3780 15056 3836
rect 14992 3776 15056 3780
rect 15072 3836 15136 3840
rect 15072 3780 15076 3836
rect 15076 3780 15132 3836
rect 15132 3780 15136 3836
rect 15072 3776 15136 3780
rect 15152 3836 15216 3840
rect 15152 3780 15156 3836
rect 15156 3780 15212 3836
rect 15212 3780 15216 3836
rect 15152 3776 15216 3780
rect 15232 3836 15296 3840
rect 15232 3780 15236 3836
rect 15236 3780 15292 3836
rect 15292 3780 15296 3836
rect 15232 3776 15296 3780
rect 18912 3836 18976 3840
rect 18912 3780 18916 3836
rect 18916 3780 18972 3836
rect 18972 3780 18976 3836
rect 18912 3776 18976 3780
rect 18992 3836 19056 3840
rect 18992 3780 18996 3836
rect 18996 3780 19052 3836
rect 19052 3780 19056 3836
rect 18992 3776 19056 3780
rect 19072 3836 19136 3840
rect 19072 3780 19076 3836
rect 19076 3780 19132 3836
rect 19132 3780 19136 3836
rect 19072 3776 19136 3780
rect 19152 3836 19216 3840
rect 19152 3780 19156 3836
rect 19156 3780 19212 3836
rect 19212 3780 19216 3836
rect 19152 3776 19216 3780
rect 19232 3836 19296 3840
rect 19232 3780 19236 3836
rect 19236 3780 19292 3836
rect 19292 3780 19296 3836
rect 19232 3776 19296 3780
rect 22912 3836 22976 3840
rect 22912 3780 22916 3836
rect 22916 3780 22972 3836
rect 22972 3780 22976 3836
rect 22912 3776 22976 3780
rect 22992 3836 23056 3840
rect 22992 3780 22996 3836
rect 22996 3780 23052 3836
rect 23052 3780 23056 3836
rect 22992 3776 23056 3780
rect 23072 3836 23136 3840
rect 23072 3780 23076 3836
rect 23076 3780 23132 3836
rect 23132 3780 23136 3836
rect 23072 3776 23136 3780
rect 23152 3836 23216 3840
rect 23152 3780 23156 3836
rect 23156 3780 23212 3836
rect 23212 3780 23216 3836
rect 23152 3776 23216 3780
rect 23232 3836 23296 3840
rect 23232 3780 23236 3836
rect 23236 3780 23292 3836
rect 23292 3780 23296 3836
rect 23232 3776 23296 3780
rect 3652 3292 3716 3296
rect 3652 3236 3656 3292
rect 3656 3236 3712 3292
rect 3712 3236 3716 3292
rect 3652 3232 3716 3236
rect 3732 3292 3796 3296
rect 3732 3236 3736 3292
rect 3736 3236 3792 3292
rect 3792 3236 3796 3292
rect 3732 3232 3796 3236
rect 3812 3292 3876 3296
rect 3812 3236 3816 3292
rect 3816 3236 3872 3292
rect 3872 3236 3876 3292
rect 3812 3232 3876 3236
rect 3892 3292 3956 3296
rect 3892 3236 3896 3292
rect 3896 3236 3952 3292
rect 3952 3236 3956 3292
rect 3892 3232 3956 3236
rect 3972 3292 4036 3296
rect 3972 3236 3976 3292
rect 3976 3236 4032 3292
rect 4032 3236 4036 3292
rect 3972 3232 4036 3236
rect 7652 3292 7716 3296
rect 7652 3236 7656 3292
rect 7656 3236 7712 3292
rect 7712 3236 7716 3292
rect 7652 3232 7716 3236
rect 7732 3292 7796 3296
rect 7732 3236 7736 3292
rect 7736 3236 7792 3292
rect 7792 3236 7796 3292
rect 7732 3232 7796 3236
rect 7812 3292 7876 3296
rect 7812 3236 7816 3292
rect 7816 3236 7872 3292
rect 7872 3236 7876 3292
rect 7812 3232 7876 3236
rect 7892 3292 7956 3296
rect 7892 3236 7896 3292
rect 7896 3236 7952 3292
rect 7952 3236 7956 3292
rect 7892 3232 7956 3236
rect 7972 3292 8036 3296
rect 7972 3236 7976 3292
rect 7976 3236 8032 3292
rect 8032 3236 8036 3292
rect 7972 3232 8036 3236
rect 11652 3292 11716 3296
rect 11652 3236 11656 3292
rect 11656 3236 11712 3292
rect 11712 3236 11716 3292
rect 11652 3232 11716 3236
rect 11732 3292 11796 3296
rect 11732 3236 11736 3292
rect 11736 3236 11792 3292
rect 11792 3236 11796 3292
rect 11732 3232 11796 3236
rect 11812 3292 11876 3296
rect 11812 3236 11816 3292
rect 11816 3236 11872 3292
rect 11872 3236 11876 3292
rect 11812 3232 11876 3236
rect 11892 3292 11956 3296
rect 11892 3236 11896 3292
rect 11896 3236 11952 3292
rect 11952 3236 11956 3292
rect 11892 3232 11956 3236
rect 11972 3292 12036 3296
rect 11972 3236 11976 3292
rect 11976 3236 12032 3292
rect 12032 3236 12036 3292
rect 11972 3232 12036 3236
rect 15652 3292 15716 3296
rect 15652 3236 15656 3292
rect 15656 3236 15712 3292
rect 15712 3236 15716 3292
rect 15652 3232 15716 3236
rect 15732 3292 15796 3296
rect 15732 3236 15736 3292
rect 15736 3236 15792 3292
rect 15792 3236 15796 3292
rect 15732 3232 15796 3236
rect 15812 3292 15876 3296
rect 15812 3236 15816 3292
rect 15816 3236 15872 3292
rect 15872 3236 15876 3292
rect 15812 3232 15876 3236
rect 15892 3292 15956 3296
rect 15892 3236 15896 3292
rect 15896 3236 15952 3292
rect 15952 3236 15956 3292
rect 15892 3232 15956 3236
rect 15972 3292 16036 3296
rect 15972 3236 15976 3292
rect 15976 3236 16032 3292
rect 16032 3236 16036 3292
rect 15972 3232 16036 3236
rect 19652 3292 19716 3296
rect 19652 3236 19656 3292
rect 19656 3236 19712 3292
rect 19712 3236 19716 3292
rect 19652 3232 19716 3236
rect 19732 3292 19796 3296
rect 19732 3236 19736 3292
rect 19736 3236 19792 3292
rect 19792 3236 19796 3292
rect 19732 3232 19796 3236
rect 19812 3292 19876 3296
rect 19812 3236 19816 3292
rect 19816 3236 19872 3292
rect 19872 3236 19876 3292
rect 19812 3232 19876 3236
rect 19892 3292 19956 3296
rect 19892 3236 19896 3292
rect 19896 3236 19952 3292
rect 19952 3236 19956 3292
rect 19892 3232 19956 3236
rect 19972 3292 20036 3296
rect 19972 3236 19976 3292
rect 19976 3236 20032 3292
rect 20032 3236 20036 3292
rect 19972 3232 20036 3236
rect 23652 3292 23716 3296
rect 23652 3236 23656 3292
rect 23656 3236 23712 3292
rect 23712 3236 23716 3292
rect 23652 3232 23716 3236
rect 23732 3292 23796 3296
rect 23732 3236 23736 3292
rect 23736 3236 23792 3292
rect 23792 3236 23796 3292
rect 23732 3232 23796 3236
rect 23812 3292 23876 3296
rect 23812 3236 23816 3292
rect 23816 3236 23872 3292
rect 23872 3236 23876 3292
rect 23812 3232 23876 3236
rect 23892 3292 23956 3296
rect 23892 3236 23896 3292
rect 23896 3236 23952 3292
rect 23952 3236 23956 3292
rect 23892 3232 23956 3236
rect 23972 3292 24036 3296
rect 23972 3236 23976 3292
rect 23976 3236 24032 3292
rect 24032 3236 24036 3292
rect 23972 3232 24036 3236
rect 2912 2748 2976 2752
rect 2912 2692 2916 2748
rect 2916 2692 2972 2748
rect 2972 2692 2976 2748
rect 2912 2688 2976 2692
rect 2992 2748 3056 2752
rect 2992 2692 2996 2748
rect 2996 2692 3052 2748
rect 3052 2692 3056 2748
rect 2992 2688 3056 2692
rect 3072 2748 3136 2752
rect 3072 2692 3076 2748
rect 3076 2692 3132 2748
rect 3132 2692 3136 2748
rect 3072 2688 3136 2692
rect 3152 2748 3216 2752
rect 3152 2692 3156 2748
rect 3156 2692 3212 2748
rect 3212 2692 3216 2748
rect 3152 2688 3216 2692
rect 3232 2748 3296 2752
rect 3232 2692 3236 2748
rect 3236 2692 3292 2748
rect 3292 2692 3296 2748
rect 3232 2688 3296 2692
rect 6912 2748 6976 2752
rect 6912 2692 6916 2748
rect 6916 2692 6972 2748
rect 6972 2692 6976 2748
rect 6912 2688 6976 2692
rect 6992 2748 7056 2752
rect 6992 2692 6996 2748
rect 6996 2692 7052 2748
rect 7052 2692 7056 2748
rect 6992 2688 7056 2692
rect 7072 2748 7136 2752
rect 7072 2692 7076 2748
rect 7076 2692 7132 2748
rect 7132 2692 7136 2748
rect 7072 2688 7136 2692
rect 7152 2748 7216 2752
rect 7152 2692 7156 2748
rect 7156 2692 7212 2748
rect 7212 2692 7216 2748
rect 7152 2688 7216 2692
rect 7232 2748 7296 2752
rect 7232 2692 7236 2748
rect 7236 2692 7292 2748
rect 7292 2692 7296 2748
rect 7232 2688 7296 2692
rect 10912 2748 10976 2752
rect 10912 2692 10916 2748
rect 10916 2692 10972 2748
rect 10972 2692 10976 2748
rect 10912 2688 10976 2692
rect 10992 2748 11056 2752
rect 10992 2692 10996 2748
rect 10996 2692 11052 2748
rect 11052 2692 11056 2748
rect 10992 2688 11056 2692
rect 11072 2748 11136 2752
rect 11072 2692 11076 2748
rect 11076 2692 11132 2748
rect 11132 2692 11136 2748
rect 11072 2688 11136 2692
rect 11152 2748 11216 2752
rect 11152 2692 11156 2748
rect 11156 2692 11212 2748
rect 11212 2692 11216 2748
rect 11152 2688 11216 2692
rect 11232 2748 11296 2752
rect 11232 2692 11236 2748
rect 11236 2692 11292 2748
rect 11292 2692 11296 2748
rect 11232 2688 11296 2692
rect 14912 2748 14976 2752
rect 14912 2692 14916 2748
rect 14916 2692 14972 2748
rect 14972 2692 14976 2748
rect 14912 2688 14976 2692
rect 14992 2748 15056 2752
rect 14992 2692 14996 2748
rect 14996 2692 15052 2748
rect 15052 2692 15056 2748
rect 14992 2688 15056 2692
rect 15072 2748 15136 2752
rect 15072 2692 15076 2748
rect 15076 2692 15132 2748
rect 15132 2692 15136 2748
rect 15072 2688 15136 2692
rect 15152 2748 15216 2752
rect 15152 2692 15156 2748
rect 15156 2692 15212 2748
rect 15212 2692 15216 2748
rect 15152 2688 15216 2692
rect 15232 2748 15296 2752
rect 15232 2692 15236 2748
rect 15236 2692 15292 2748
rect 15292 2692 15296 2748
rect 15232 2688 15296 2692
rect 18912 2748 18976 2752
rect 18912 2692 18916 2748
rect 18916 2692 18972 2748
rect 18972 2692 18976 2748
rect 18912 2688 18976 2692
rect 18992 2748 19056 2752
rect 18992 2692 18996 2748
rect 18996 2692 19052 2748
rect 19052 2692 19056 2748
rect 18992 2688 19056 2692
rect 19072 2748 19136 2752
rect 19072 2692 19076 2748
rect 19076 2692 19132 2748
rect 19132 2692 19136 2748
rect 19072 2688 19136 2692
rect 19152 2748 19216 2752
rect 19152 2692 19156 2748
rect 19156 2692 19212 2748
rect 19212 2692 19216 2748
rect 19152 2688 19216 2692
rect 19232 2748 19296 2752
rect 19232 2692 19236 2748
rect 19236 2692 19292 2748
rect 19292 2692 19296 2748
rect 19232 2688 19296 2692
rect 22912 2748 22976 2752
rect 22912 2692 22916 2748
rect 22916 2692 22972 2748
rect 22972 2692 22976 2748
rect 22912 2688 22976 2692
rect 22992 2748 23056 2752
rect 22992 2692 22996 2748
rect 22996 2692 23052 2748
rect 23052 2692 23056 2748
rect 22992 2688 23056 2692
rect 23072 2748 23136 2752
rect 23072 2692 23076 2748
rect 23076 2692 23132 2748
rect 23132 2692 23136 2748
rect 23072 2688 23136 2692
rect 23152 2748 23216 2752
rect 23152 2692 23156 2748
rect 23156 2692 23212 2748
rect 23212 2692 23216 2748
rect 23152 2688 23216 2692
rect 23232 2748 23296 2752
rect 23232 2692 23236 2748
rect 23236 2692 23292 2748
rect 23292 2692 23296 2748
rect 23232 2688 23296 2692
rect 3652 2204 3716 2208
rect 3652 2148 3656 2204
rect 3656 2148 3712 2204
rect 3712 2148 3716 2204
rect 3652 2144 3716 2148
rect 3732 2204 3796 2208
rect 3732 2148 3736 2204
rect 3736 2148 3792 2204
rect 3792 2148 3796 2204
rect 3732 2144 3796 2148
rect 3812 2204 3876 2208
rect 3812 2148 3816 2204
rect 3816 2148 3872 2204
rect 3872 2148 3876 2204
rect 3812 2144 3876 2148
rect 3892 2204 3956 2208
rect 3892 2148 3896 2204
rect 3896 2148 3952 2204
rect 3952 2148 3956 2204
rect 3892 2144 3956 2148
rect 3972 2204 4036 2208
rect 3972 2148 3976 2204
rect 3976 2148 4032 2204
rect 4032 2148 4036 2204
rect 3972 2144 4036 2148
rect 7652 2204 7716 2208
rect 7652 2148 7656 2204
rect 7656 2148 7712 2204
rect 7712 2148 7716 2204
rect 7652 2144 7716 2148
rect 7732 2204 7796 2208
rect 7732 2148 7736 2204
rect 7736 2148 7792 2204
rect 7792 2148 7796 2204
rect 7732 2144 7796 2148
rect 7812 2204 7876 2208
rect 7812 2148 7816 2204
rect 7816 2148 7872 2204
rect 7872 2148 7876 2204
rect 7812 2144 7876 2148
rect 7892 2204 7956 2208
rect 7892 2148 7896 2204
rect 7896 2148 7952 2204
rect 7952 2148 7956 2204
rect 7892 2144 7956 2148
rect 7972 2204 8036 2208
rect 7972 2148 7976 2204
rect 7976 2148 8032 2204
rect 8032 2148 8036 2204
rect 7972 2144 8036 2148
rect 11652 2204 11716 2208
rect 11652 2148 11656 2204
rect 11656 2148 11712 2204
rect 11712 2148 11716 2204
rect 11652 2144 11716 2148
rect 11732 2204 11796 2208
rect 11732 2148 11736 2204
rect 11736 2148 11792 2204
rect 11792 2148 11796 2204
rect 11732 2144 11796 2148
rect 11812 2204 11876 2208
rect 11812 2148 11816 2204
rect 11816 2148 11872 2204
rect 11872 2148 11876 2204
rect 11812 2144 11876 2148
rect 11892 2204 11956 2208
rect 11892 2148 11896 2204
rect 11896 2148 11952 2204
rect 11952 2148 11956 2204
rect 11892 2144 11956 2148
rect 11972 2204 12036 2208
rect 11972 2148 11976 2204
rect 11976 2148 12032 2204
rect 12032 2148 12036 2204
rect 11972 2144 12036 2148
rect 15652 2204 15716 2208
rect 15652 2148 15656 2204
rect 15656 2148 15712 2204
rect 15712 2148 15716 2204
rect 15652 2144 15716 2148
rect 15732 2204 15796 2208
rect 15732 2148 15736 2204
rect 15736 2148 15792 2204
rect 15792 2148 15796 2204
rect 15732 2144 15796 2148
rect 15812 2204 15876 2208
rect 15812 2148 15816 2204
rect 15816 2148 15872 2204
rect 15872 2148 15876 2204
rect 15812 2144 15876 2148
rect 15892 2204 15956 2208
rect 15892 2148 15896 2204
rect 15896 2148 15952 2204
rect 15952 2148 15956 2204
rect 15892 2144 15956 2148
rect 15972 2204 16036 2208
rect 15972 2148 15976 2204
rect 15976 2148 16032 2204
rect 16032 2148 16036 2204
rect 15972 2144 16036 2148
rect 19652 2204 19716 2208
rect 19652 2148 19656 2204
rect 19656 2148 19712 2204
rect 19712 2148 19716 2204
rect 19652 2144 19716 2148
rect 19732 2204 19796 2208
rect 19732 2148 19736 2204
rect 19736 2148 19792 2204
rect 19792 2148 19796 2204
rect 19732 2144 19796 2148
rect 19812 2204 19876 2208
rect 19812 2148 19816 2204
rect 19816 2148 19872 2204
rect 19872 2148 19876 2204
rect 19812 2144 19876 2148
rect 19892 2204 19956 2208
rect 19892 2148 19896 2204
rect 19896 2148 19952 2204
rect 19952 2148 19956 2204
rect 19892 2144 19956 2148
rect 19972 2204 20036 2208
rect 19972 2148 19976 2204
rect 19976 2148 20032 2204
rect 20032 2148 20036 2204
rect 19972 2144 20036 2148
rect 23652 2204 23716 2208
rect 23652 2148 23656 2204
rect 23656 2148 23712 2204
rect 23712 2148 23716 2204
rect 23652 2144 23716 2148
rect 23732 2204 23796 2208
rect 23732 2148 23736 2204
rect 23736 2148 23792 2204
rect 23792 2148 23796 2204
rect 23732 2144 23796 2148
rect 23812 2204 23876 2208
rect 23812 2148 23816 2204
rect 23816 2148 23872 2204
rect 23872 2148 23876 2204
rect 23812 2144 23876 2148
rect 23892 2204 23956 2208
rect 23892 2148 23896 2204
rect 23896 2148 23952 2204
rect 23952 2148 23956 2204
rect 23892 2144 23956 2148
rect 23972 2204 24036 2208
rect 23972 2148 23976 2204
rect 23976 2148 24032 2204
rect 24032 2148 24036 2204
rect 23972 2144 24036 2148
<< metal4 >>
rect 2904 27776 3304 27792
rect 2904 27712 2912 27776
rect 2976 27712 2992 27776
rect 3056 27712 3072 27776
rect 3136 27712 3152 27776
rect 3216 27712 3232 27776
rect 3296 27712 3304 27776
rect 2904 26688 3304 27712
rect 2904 26624 2912 26688
rect 2976 26624 2992 26688
rect 3056 26624 3072 26688
rect 3136 26624 3152 26688
rect 3216 26624 3232 26688
rect 3296 26624 3304 26688
rect 2904 25600 3304 26624
rect 2904 25536 2912 25600
rect 2976 25536 2992 25600
rect 3056 25536 3072 25600
rect 3136 25536 3152 25600
rect 3216 25536 3232 25600
rect 3296 25536 3304 25600
rect 2904 24512 3304 25536
rect 2904 24448 2912 24512
rect 2976 24448 2992 24512
rect 3056 24448 3072 24512
rect 3136 24448 3152 24512
rect 3216 24448 3232 24512
rect 3296 24448 3304 24512
rect 2904 24294 3304 24448
rect 2904 24058 2986 24294
rect 3222 24058 3304 24294
rect 2904 23424 3304 24058
rect 2904 23360 2912 23424
rect 2976 23360 2992 23424
rect 3056 23360 3072 23424
rect 3136 23360 3152 23424
rect 3216 23360 3232 23424
rect 3296 23360 3304 23424
rect 2904 22336 3304 23360
rect 2904 22272 2912 22336
rect 2976 22272 2992 22336
rect 3056 22272 3072 22336
rect 3136 22272 3152 22336
rect 3216 22272 3232 22336
rect 3296 22272 3304 22336
rect 2904 21248 3304 22272
rect 2904 21184 2912 21248
rect 2976 21184 2992 21248
rect 3056 21184 3072 21248
rect 3136 21184 3152 21248
rect 3216 21184 3232 21248
rect 3296 21184 3304 21248
rect 2904 20294 3304 21184
rect 2904 20160 2986 20294
rect 3222 20160 3304 20294
rect 2904 20096 2912 20160
rect 2976 20096 2986 20160
rect 3222 20096 3232 20160
rect 3296 20096 3304 20160
rect 2904 20058 2986 20096
rect 3222 20058 3304 20096
rect 2904 19072 3304 20058
rect 2904 19008 2912 19072
rect 2976 19008 2992 19072
rect 3056 19008 3072 19072
rect 3136 19008 3152 19072
rect 3216 19008 3232 19072
rect 3296 19008 3304 19072
rect 2904 17984 3304 19008
rect 2904 17920 2912 17984
rect 2976 17920 2992 17984
rect 3056 17920 3072 17984
rect 3136 17920 3152 17984
rect 3216 17920 3232 17984
rect 3296 17920 3304 17984
rect 2904 16896 3304 17920
rect 2904 16832 2912 16896
rect 2976 16832 2992 16896
rect 3056 16832 3072 16896
rect 3136 16832 3152 16896
rect 3216 16832 3232 16896
rect 3296 16832 3304 16896
rect 2904 16294 3304 16832
rect 2904 16058 2986 16294
rect 3222 16058 3304 16294
rect 2904 15808 3304 16058
rect 2904 15744 2912 15808
rect 2976 15744 2992 15808
rect 3056 15744 3072 15808
rect 3136 15744 3152 15808
rect 3216 15744 3232 15808
rect 3296 15744 3304 15808
rect 2904 14720 3304 15744
rect 2904 14656 2912 14720
rect 2976 14656 2992 14720
rect 3056 14656 3072 14720
rect 3136 14656 3152 14720
rect 3216 14656 3232 14720
rect 3296 14656 3304 14720
rect 2904 13632 3304 14656
rect 2904 13568 2912 13632
rect 2976 13568 2992 13632
rect 3056 13568 3072 13632
rect 3136 13568 3152 13632
rect 3216 13568 3232 13632
rect 3296 13568 3304 13632
rect 2904 12544 3304 13568
rect 2904 12480 2912 12544
rect 2976 12480 2992 12544
rect 3056 12480 3072 12544
rect 3136 12480 3152 12544
rect 3216 12480 3232 12544
rect 3296 12480 3304 12544
rect 2904 12294 3304 12480
rect 2904 12058 2986 12294
rect 3222 12058 3304 12294
rect 2904 11456 3304 12058
rect 2904 11392 2912 11456
rect 2976 11392 2992 11456
rect 3056 11392 3072 11456
rect 3136 11392 3152 11456
rect 3216 11392 3232 11456
rect 3296 11392 3304 11456
rect 2904 10368 3304 11392
rect 2904 10304 2912 10368
rect 2976 10304 2992 10368
rect 3056 10304 3072 10368
rect 3136 10304 3152 10368
rect 3216 10304 3232 10368
rect 3296 10304 3304 10368
rect 2904 9280 3304 10304
rect 2904 9216 2912 9280
rect 2976 9216 2992 9280
rect 3056 9216 3072 9280
rect 3136 9216 3152 9280
rect 3216 9216 3232 9280
rect 3296 9216 3304 9280
rect 2904 8294 3304 9216
rect 2904 8192 2986 8294
rect 3222 8192 3304 8294
rect 2904 8128 2912 8192
rect 2976 8128 2986 8192
rect 3222 8128 3232 8192
rect 3296 8128 3304 8192
rect 2904 8058 2986 8128
rect 3222 8058 3304 8128
rect 2904 7104 3304 8058
rect 2904 7040 2912 7104
rect 2976 7040 2992 7104
rect 3056 7040 3072 7104
rect 3136 7040 3152 7104
rect 3216 7040 3232 7104
rect 3296 7040 3304 7104
rect 2904 6016 3304 7040
rect 2904 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3072 6016
rect 3136 5952 3152 6016
rect 3216 5952 3232 6016
rect 3296 5952 3304 6016
rect 2904 4928 3304 5952
rect 2904 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3072 4928
rect 3136 4864 3152 4928
rect 3216 4864 3232 4928
rect 3296 4864 3304 4928
rect 2904 4294 3304 4864
rect 2904 4058 2986 4294
rect 3222 4058 3304 4294
rect 2904 3840 3304 4058
rect 2904 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3072 3840
rect 3136 3776 3152 3840
rect 3216 3776 3232 3840
rect 3296 3776 3304 3840
rect 2904 2752 3304 3776
rect 2904 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3072 2752
rect 3136 2688 3152 2752
rect 3216 2688 3232 2752
rect 3296 2688 3304 2752
rect 2904 2128 3304 2688
rect 3644 27232 4044 27792
rect 3644 27168 3652 27232
rect 3716 27168 3732 27232
rect 3796 27168 3812 27232
rect 3876 27168 3892 27232
rect 3956 27168 3972 27232
rect 4036 27168 4044 27232
rect 3644 26144 4044 27168
rect 3644 26080 3652 26144
rect 3716 26080 3732 26144
rect 3796 26080 3812 26144
rect 3876 26080 3892 26144
rect 3956 26080 3972 26144
rect 4036 26080 4044 26144
rect 3644 25056 4044 26080
rect 3644 24992 3652 25056
rect 3716 25034 3732 25056
rect 3796 25034 3812 25056
rect 3876 25034 3892 25056
rect 3956 25034 3972 25056
rect 3716 24992 3726 25034
rect 3962 24992 3972 25034
rect 4036 24992 4044 25056
rect 3644 24798 3726 24992
rect 3962 24798 4044 24992
rect 3644 23968 4044 24798
rect 3644 23904 3652 23968
rect 3716 23904 3732 23968
rect 3796 23904 3812 23968
rect 3876 23904 3892 23968
rect 3956 23904 3972 23968
rect 4036 23904 4044 23968
rect 3644 22880 4044 23904
rect 3644 22816 3652 22880
rect 3716 22816 3732 22880
rect 3796 22816 3812 22880
rect 3876 22816 3892 22880
rect 3956 22816 3972 22880
rect 4036 22816 4044 22880
rect 3644 21792 4044 22816
rect 6904 27776 7304 27792
rect 6904 27712 6912 27776
rect 6976 27712 6992 27776
rect 7056 27712 7072 27776
rect 7136 27712 7152 27776
rect 7216 27712 7232 27776
rect 7296 27712 7304 27776
rect 6904 26688 7304 27712
rect 6904 26624 6912 26688
rect 6976 26624 6992 26688
rect 7056 26624 7072 26688
rect 7136 26624 7152 26688
rect 7216 26624 7232 26688
rect 7296 26624 7304 26688
rect 6904 25600 7304 26624
rect 6904 25536 6912 25600
rect 6976 25536 6992 25600
rect 7056 25536 7072 25600
rect 7136 25536 7152 25600
rect 7216 25536 7232 25600
rect 7296 25536 7304 25600
rect 6904 24512 7304 25536
rect 6904 24448 6912 24512
rect 6976 24448 6992 24512
rect 7056 24448 7072 24512
rect 7136 24448 7152 24512
rect 7216 24448 7232 24512
rect 7296 24448 7304 24512
rect 6904 24294 7304 24448
rect 6904 24058 6986 24294
rect 7222 24058 7304 24294
rect 6904 23424 7304 24058
rect 6904 23360 6912 23424
rect 6976 23360 6992 23424
rect 7056 23360 7072 23424
rect 7136 23360 7152 23424
rect 7216 23360 7232 23424
rect 7296 23360 7304 23424
rect 6904 22336 7304 23360
rect 6904 22272 6912 22336
rect 6976 22272 6992 22336
rect 7056 22272 7072 22336
rect 7136 22272 7152 22336
rect 7216 22272 7232 22336
rect 7296 22272 7304 22336
rect 5395 22132 5461 22133
rect 5395 22068 5396 22132
rect 5460 22068 5461 22132
rect 5395 22067 5461 22068
rect 3644 21728 3652 21792
rect 3716 21728 3732 21792
rect 3796 21728 3812 21792
rect 3876 21728 3892 21792
rect 3956 21728 3972 21792
rect 4036 21728 4044 21792
rect 3644 21034 4044 21728
rect 3644 20798 3726 21034
rect 3962 20798 4044 21034
rect 3644 20704 4044 20798
rect 3644 20640 3652 20704
rect 3716 20640 3732 20704
rect 3796 20640 3812 20704
rect 3876 20640 3892 20704
rect 3956 20640 3972 20704
rect 4036 20640 4044 20704
rect 3644 19616 4044 20640
rect 3644 19552 3652 19616
rect 3716 19552 3732 19616
rect 3796 19552 3812 19616
rect 3876 19552 3892 19616
rect 3956 19552 3972 19616
rect 4036 19552 4044 19616
rect 3644 18528 4044 19552
rect 5211 19412 5277 19413
rect 5211 19348 5212 19412
rect 5276 19348 5277 19412
rect 5211 19347 5277 19348
rect 3644 18464 3652 18528
rect 3716 18464 3732 18528
rect 3796 18464 3812 18528
rect 3876 18464 3892 18528
rect 3956 18464 3972 18528
rect 4036 18464 4044 18528
rect 3644 17440 4044 18464
rect 3644 17376 3652 17440
rect 3716 17376 3732 17440
rect 3796 17376 3812 17440
rect 3876 17376 3892 17440
rect 3956 17376 3972 17440
rect 4036 17376 4044 17440
rect 3644 17034 4044 17376
rect 3644 16798 3726 17034
rect 3962 16798 4044 17034
rect 3644 16352 4044 16798
rect 3644 16288 3652 16352
rect 3716 16288 3732 16352
rect 3796 16288 3812 16352
rect 3876 16288 3892 16352
rect 3956 16288 3972 16352
rect 4036 16288 4044 16352
rect 3644 15264 4044 16288
rect 3644 15200 3652 15264
rect 3716 15200 3732 15264
rect 3796 15200 3812 15264
rect 3876 15200 3892 15264
rect 3956 15200 3972 15264
rect 4036 15200 4044 15264
rect 3644 14176 4044 15200
rect 3644 14112 3652 14176
rect 3716 14112 3732 14176
rect 3796 14112 3812 14176
rect 3876 14112 3892 14176
rect 3956 14112 3972 14176
rect 4036 14112 4044 14176
rect 3644 13088 4044 14112
rect 3644 13024 3652 13088
rect 3716 13034 3732 13088
rect 3796 13034 3812 13088
rect 3876 13034 3892 13088
rect 3956 13034 3972 13088
rect 3716 13024 3726 13034
rect 3962 13024 3972 13034
rect 4036 13024 4044 13088
rect 3644 12798 3726 13024
rect 3962 12798 4044 13024
rect 5214 12885 5274 19347
rect 5211 12884 5277 12885
rect 5211 12820 5212 12884
rect 5276 12820 5277 12884
rect 5211 12819 5277 12820
rect 3644 12000 4044 12798
rect 3644 11936 3652 12000
rect 3716 11936 3732 12000
rect 3796 11936 3812 12000
rect 3876 11936 3892 12000
rect 3956 11936 3972 12000
rect 4036 11936 4044 12000
rect 3644 10912 4044 11936
rect 3644 10848 3652 10912
rect 3716 10848 3732 10912
rect 3796 10848 3812 10912
rect 3876 10848 3892 10912
rect 3956 10848 3972 10912
rect 4036 10848 4044 10912
rect 3644 9824 4044 10848
rect 3644 9760 3652 9824
rect 3716 9760 3732 9824
rect 3796 9760 3812 9824
rect 3876 9760 3892 9824
rect 3956 9760 3972 9824
rect 4036 9760 4044 9824
rect 3644 9034 4044 9760
rect 3644 8798 3726 9034
rect 3962 8798 4044 9034
rect 3644 8736 4044 8798
rect 3644 8672 3652 8736
rect 3716 8672 3732 8736
rect 3796 8672 3812 8736
rect 3876 8672 3892 8736
rect 3956 8672 3972 8736
rect 4036 8672 4044 8736
rect 3644 7648 4044 8672
rect 3644 7584 3652 7648
rect 3716 7584 3732 7648
rect 3796 7584 3812 7648
rect 3876 7584 3892 7648
rect 3956 7584 3972 7648
rect 4036 7584 4044 7648
rect 3644 6560 4044 7584
rect 5214 7037 5274 12819
rect 5398 11797 5458 22067
rect 6904 21248 7304 22272
rect 6904 21184 6912 21248
rect 6976 21184 6992 21248
rect 7056 21184 7072 21248
rect 7136 21184 7152 21248
rect 7216 21184 7232 21248
rect 7296 21184 7304 21248
rect 6904 20294 7304 21184
rect 6904 20160 6986 20294
rect 7222 20160 7304 20294
rect 6904 20096 6912 20160
rect 6976 20096 6986 20160
rect 7222 20096 7232 20160
rect 7296 20096 7304 20160
rect 6904 20058 6986 20096
rect 7222 20058 7304 20096
rect 6904 19072 7304 20058
rect 6904 19008 6912 19072
rect 6976 19008 6992 19072
rect 7056 19008 7072 19072
rect 7136 19008 7152 19072
rect 7216 19008 7232 19072
rect 7296 19008 7304 19072
rect 6904 17984 7304 19008
rect 6904 17920 6912 17984
rect 6976 17920 6992 17984
rect 7056 17920 7072 17984
rect 7136 17920 7152 17984
rect 7216 17920 7232 17984
rect 7296 17920 7304 17984
rect 6904 16896 7304 17920
rect 6904 16832 6912 16896
rect 6976 16832 6992 16896
rect 7056 16832 7072 16896
rect 7136 16832 7152 16896
rect 7216 16832 7232 16896
rect 7296 16832 7304 16896
rect 6904 16294 7304 16832
rect 6904 16058 6986 16294
rect 7222 16058 7304 16294
rect 6904 15808 7304 16058
rect 6904 15744 6912 15808
rect 6976 15744 6992 15808
rect 7056 15744 7072 15808
rect 7136 15744 7152 15808
rect 7216 15744 7232 15808
rect 7296 15744 7304 15808
rect 6904 14720 7304 15744
rect 6904 14656 6912 14720
rect 6976 14656 6992 14720
rect 7056 14656 7072 14720
rect 7136 14656 7152 14720
rect 7216 14656 7232 14720
rect 7296 14656 7304 14720
rect 6904 13632 7304 14656
rect 6904 13568 6912 13632
rect 6976 13568 6992 13632
rect 7056 13568 7072 13632
rect 7136 13568 7152 13632
rect 7216 13568 7232 13632
rect 7296 13568 7304 13632
rect 6904 12544 7304 13568
rect 6904 12480 6912 12544
rect 6976 12480 6992 12544
rect 7056 12480 7072 12544
rect 7136 12480 7152 12544
rect 7216 12480 7232 12544
rect 7296 12480 7304 12544
rect 6904 12294 7304 12480
rect 6904 12058 6986 12294
rect 7222 12058 7304 12294
rect 5395 11796 5461 11797
rect 5395 11732 5396 11796
rect 5460 11732 5461 11796
rect 5395 11731 5461 11732
rect 6904 11456 7304 12058
rect 6904 11392 6912 11456
rect 6976 11392 6992 11456
rect 7056 11392 7072 11456
rect 7136 11392 7152 11456
rect 7216 11392 7232 11456
rect 7296 11392 7304 11456
rect 6904 10368 7304 11392
rect 6904 10304 6912 10368
rect 6976 10304 6992 10368
rect 7056 10304 7072 10368
rect 7136 10304 7152 10368
rect 7216 10304 7232 10368
rect 7296 10304 7304 10368
rect 6904 9280 7304 10304
rect 6904 9216 6912 9280
rect 6976 9216 6992 9280
rect 7056 9216 7072 9280
rect 7136 9216 7152 9280
rect 7216 9216 7232 9280
rect 7296 9216 7304 9280
rect 6904 8294 7304 9216
rect 6904 8192 6986 8294
rect 7222 8192 7304 8294
rect 6904 8128 6912 8192
rect 6976 8128 6986 8192
rect 7222 8128 7232 8192
rect 7296 8128 7304 8192
rect 6904 8058 6986 8128
rect 7222 8058 7304 8128
rect 6904 7104 7304 8058
rect 6904 7040 6912 7104
rect 6976 7040 6992 7104
rect 7056 7040 7072 7104
rect 7136 7040 7152 7104
rect 7216 7040 7232 7104
rect 7296 7040 7304 7104
rect 5211 7036 5277 7037
rect 5211 6972 5212 7036
rect 5276 6972 5277 7036
rect 5211 6971 5277 6972
rect 3644 6496 3652 6560
rect 3716 6496 3732 6560
rect 3796 6496 3812 6560
rect 3876 6496 3892 6560
rect 3956 6496 3972 6560
rect 4036 6496 4044 6560
rect 3644 5472 4044 6496
rect 3644 5408 3652 5472
rect 3716 5408 3732 5472
rect 3796 5408 3812 5472
rect 3876 5408 3892 5472
rect 3956 5408 3972 5472
rect 4036 5408 4044 5472
rect 3644 5034 4044 5408
rect 3644 4798 3726 5034
rect 3962 4798 4044 5034
rect 3644 4384 4044 4798
rect 3644 4320 3652 4384
rect 3716 4320 3732 4384
rect 3796 4320 3812 4384
rect 3876 4320 3892 4384
rect 3956 4320 3972 4384
rect 4036 4320 4044 4384
rect 3644 3296 4044 4320
rect 3644 3232 3652 3296
rect 3716 3232 3732 3296
rect 3796 3232 3812 3296
rect 3876 3232 3892 3296
rect 3956 3232 3972 3296
rect 4036 3232 4044 3296
rect 3644 2208 4044 3232
rect 3644 2144 3652 2208
rect 3716 2144 3732 2208
rect 3796 2144 3812 2208
rect 3876 2144 3892 2208
rect 3956 2144 3972 2208
rect 4036 2144 4044 2208
rect 3644 2128 4044 2144
rect 6904 6016 7304 7040
rect 6904 5952 6912 6016
rect 6976 5952 6992 6016
rect 7056 5952 7072 6016
rect 7136 5952 7152 6016
rect 7216 5952 7232 6016
rect 7296 5952 7304 6016
rect 6904 4928 7304 5952
rect 6904 4864 6912 4928
rect 6976 4864 6992 4928
rect 7056 4864 7072 4928
rect 7136 4864 7152 4928
rect 7216 4864 7232 4928
rect 7296 4864 7304 4928
rect 6904 4294 7304 4864
rect 6904 4058 6986 4294
rect 7222 4058 7304 4294
rect 6904 3840 7304 4058
rect 6904 3776 6912 3840
rect 6976 3776 6992 3840
rect 7056 3776 7072 3840
rect 7136 3776 7152 3840
rect 7216 3776 7232 3840
rect 7296 3776 7304 3840
rect 6904 2752 7304 3776
rect 6904 2688 6912 2752
rect 6976 2688 6992 2752
rect 7056 2688 7072 2752
rect 7136 2688 7152 2752
rect 7216 2688 7232 2752
rect 7296 2688 7304 2752
rect 6904 2128 7304 2688
rect 7644 27232 8044 27792
rect 7644 27168 7652 27232
rect 7716 27168 7732 27232
rect 7796 27168 7812 27232
rect 7876 27168 7892 27232
rect 7956 27168 7972 27232
rect 8036 27168 8044 27232
rect 7644 26144 8044 27168
rect 10904 27776 11304 27792
rect 10904 27712 10912 27776
rect 10976 27712 10992 27776
rect 11056 27712 11072 27776
rect 11136 27712 11152 27776
rect 11216 27712 11232 27776
rect 11296 27712 11304 27776
rect 10179 26892 10245 26893
rect 10179 26828 10180 26892
rect 10244 26828 10245 26892
rect 10179 26827 10245 26828
rect 7644 26080 7652 26144
rect 7716 26080 7732 26144
rect 7796 26080 7812 26144
rect 7876 26080 7892 26144
rect 7956 26080 7972 26144
rect 8036 26080 8044 26144
rect 7644 25056 8044 26080
rect 7644 24992 7652 25056
rect 7716 25034 7732 25056
rect 7796 25034 7812 25056
rect 7876 25034 7892 25056
rect 7956 25034 7972 25056
rect 7716 24992 7726 25034
rect 7962 24992 7972 25034
rect 8036 24992 8044 25056
rect 7644 24798 7726 24992
rect 7962 24798 8044 24992
rect 7644 23968 8044 24798
rect 7644 23904 7652 23968
rect 7716 23904 7732 23968
rect 7796 23904 7812 23968
rect 7876 23904 7892 23968
rect 7956 23904 7972 23968
rect 8036 23904 8044 23968
rect 7644 22880 8044 23904
rect 7644 22816 7652 22880
rect 7716 22816 7732 22880
rect 7796 22816 7812 22880
rect 7876 22816 7892 22880
rect 7956 22816 7972 22880
rect 8036 22816 8044 22880
rect 7644 21792 8044 22816
rect 7644 21728 7652 21792
rect 7716 21728 7732 21792
rect 7796 21728 7812 21792
rect 7876 21728 7892 21792
rect 7956 21728 7972 21792
rect 8036 21728 8044 21792
rect 7644 21034 8044 21728
rect 7644 20798 7726 21034
rect 7962 20798 8044 21034
rect 7644 20704 8044 20798
rect 7644 20640 7652 20704
rect 7716 20640 7732 20704
rect 7796 20640 7812 20704
rect 7876 20640 7892 20704
rect 7956 20640 7972 20704
rect 8036 20640 8044 20704
rect 7644 19616 8044 20640
rect 7644 19552 7652 19616
rect 7716 19552 7732 19616
rect 7796 19552 7812 19616
rect 7876 19552 7892 19616
rect 7956 19552 7972 19616
rect 8036 19552 8044 19616
rect 7644 18528 8044 19552
rect 9995 19276 10061 19277
rect 9995 19212 9996 19276
rect 10060 19212 10061 19276
rect 9995 19211 10061 19212
rect 7644 18464 7652 18528
rect 7716 18464 7732 18528
rect 7796 18464 7812 18528
rect 7876 18464 7892 18528
rect 7956 18464 7972 18528
rect 8036 18464 8044 18528
rect 7644 17440 8044 18464
rect 7644 17376 7652 17440
rect 7716 17376 7732 17440
rect 7796 17376 7812 17440
rect 7876 17376 7892 17440
rect 7956 17376 7972 17440
rect 8036 17376 8044 17440
rect 7644 17034 8044 17376
rect 7644 16798 7726 17034
rect 7962 16798 8044 17034
rect 7644 16352 8044 16798
rect 7644 16288 7652 16352
rect 7716 16288 7732 16352
rect 7796 16288 7812 16352
rect 7876 16288 7892 16352
rect 7956 16288 7972 16352
rect 8036 16288 8044 16352
rect 7644 15264 8044 16288
rect 7644 15200 7652 15264
rect 7716 15200 7732 15264
rect 7796 15200 7812 15264
rect 7876 15200 7892 15264
rect 7956 15200 7972 15264
rect 8036 15200 8044 15264
rect 7644 14176 8044 15200
rect 7644 14112 7652 14176
rect 7716 14112 7732 14176
rect 7796 14112 7812 14176
rect 7876 14112 7892 14176
rect 7956 14112 7972 14176
rect 8036 14112 8044 14176
rect 7644 13088 8044 14112
rect 7644 13024 7652 13088
rect 7716 13034 7732 13088
rect 7796 13034 7812 13088
rect 7876 13034 7892 13088
rect 7956 13034 7972 13088
rect 7716 13024 7726 13034
rect 7962 13024 7972 13034
rect 8036 13024 8044 13088
rect 7644 12798 7726 13024
rect 7962 12798 8044 13024
rect 7644 12000 8044 12798
rect 7644 11936 7652 12000
rect 7716 11936 7732 12000
rect 7796 11936 7812 12000
rect 7876 11936 7892 12000
rect 7956 11936 7972 12000
rect 8036 11936 8044 12000
rect 7644 10912 8044 11936
rect 9998 11661 10058 19211
rect 9995 11660 10061 11661
rect 9995 11596 9996 11660
rect 10060 11596 10061 11660
rect 9995 11595 10061 11596
rect 7644 10848 7652 10912
rect 7716 10848 7732 10912
rect 7796 10848 7812 10912
rect 7876 10848 7892 10912
rect 7956 10848 7972 10912
rect 8036 10848 8044 10912
rect 7644 9824 8044 10848
rect 10182 10845 10242 26827
rect 10904 26688 11304 27712
rect 10904 26624 10912 26688
rect 10976 26624 10992 26688
rect 11056 26624 11072 26688
rect 11136 26624 11152 26688
rect 11216 26624 11232 26688
rect 11296 26624 11304 26688
rect 10904 25600 11304 26624
rect 10904 25536 10912 25600
rect 10976 25536 10992 25600
rect 11056 25536 11072 25600
rect 11136 25536 11152 25600
rect 11216 25536 11232 25600
rect 11296 25536 11304 25600
rect 10904 24512 11304 25536
rect 10904 24448 10912 24512
rect 10976 24448 10992 24512
rect 11056 24448 11072 24512
rect 11136 24448 11152 24512
rect 11216 24448 11232 24512
rect 11296 24448 11304 24512
rect 10904 24294 11304 24448
rect 10904 24058 10986 24294
rect 11222 24058 11304 24294
rect 10904 23424 11304 24058
rect 10904 23360 10912 23424
rect 10976 23360 10992 23424
rect 11056 23360 11072 23424
rect 11136 23360 11152 23424
rect 11216 23360 11232 23424
rect 11296 23360 11304 23424
rect 10904 22336 11304 23360
rect 10904 22272 10912 22336
rect 10976 22272 10992 22336
rect 11056 22272 11072 22336
rect 11136 22272 11152 22336
rect 11216 22272 11232 22336
rect 11296 22272 11304 22336
rect 10904 21248 11304 22272
rect 10904 21184 10912 21248
rect 10976 21184 10992 21248
rect 11056 21184 11072 21248
rect 11136 21184 11152 21248
rect 11216 21184 11232 21248
rect 11296 21184 11304 21248
rect 10904 20294 11304 21184
rect 10904 20160 10986 20294
rect 11222 20160 11304 20294
rect 10904 20096 10912 20160
rect 10976 20096 10986 20160
rect 11222 20096 11232 20160
rect 11296 20096 11304 20160
rect 10904 20058 10986 20096
rect 11222 20058 11304 20096
rect 10904 19072 11304 20058
rect 10904 19008 10912 19072
rect 10976 19008 10992 19072
rect 11056 19008 11072 19072
rect 11136 19008 11152 19072
rect 11216 19008 11232 19072
rect 11296 19008 11304 19072
rect 10904 17984 11304 19008
rect 10904 17920 10912 17984
rect 10976 17920 10992 17984
rect 11056 17920 11072 17984
rect 11136 17920 11152 17984
rect 11216 17920 11232 17984
rect 11296 17920 11304 17984
rect 10904 16896 11304 17920
rect 10904 16832 10912 16896
rect 10976 16832 10992 16896
rect 11056 16832 11072 16896
rect 11136 16832 11152 16896
rect 11216 16832 11232 16896
rect 11296 16832 11304 16896
rect 10904 16294 11304 16832
rect 10904 16058 10986 16294
rect 11222 16058 11304 16294
rect 10904 15808 11304 16058
rect 10904 15744 10912 15808
rect 10976 15744 10992 15808
rect 11056 15744 11072 15808
rect 11136 15744 11152 15808
rect 11216 15744 11232 15808
rect 11296 15744 11304 15808
rect 10904 14720 11304 15744
rect 10904 14656 10912 14720
rect 10976 14656 10992 14720
rect 11056 14656 11072 14720
rect 11136 14656 11152 14720
rect 11216 14656 11232 14720
rect 11296 14656 11304 14720
rect 10904 13632 11304 14656
rect 10904 13568 10912 13632
rect 10976 13568 10992 13632
rect 11056 13568 11072 13632
rect 11136 13568 11152 13632
rect 11216 13568 11232 13632
rect 11296 13568 11304 13632
rect 10904 12544 11304 13568
rect 10904 12480 10912 12544
rect 10976 12480 10992 12544
rect 11056 12480 11072 12544
rect 11136 12480 11152 12544
rect 11216 12480 11232 12544
rect 11296 12480 11304 12544
rect 10904 12294 11304 12480
rect 10904 12058 10986 12294
rect 11222 12058 11304 12294
rect 10904 11456 11304 12058
rect 10904 11392 10912 11456
rect 10976 11392 10992 11456
rect 11056 11392 11072 11456
rect 11136 11392 11152 11456
rect 11216 11392 11232 11456
rect 11296 11392 11304 11456
rect 10179 10844 10245 10845
rect 10179 10780 10180 10844
rect 10244 10780 10245 10844
rect 10179 10779 10245 10780
rect 7644 9760 7652 9824
rect 7716 9760 7732 9824
rect 7796 9760 7812 9824
rect 7876 9760 7892 9824
rect 7956 9760 7972 9824
rect 8036 9760 8044 9824
rect 7644 9034 8044 9760
rect 7644 8798 7726 9034
rect 7962 8798 8044 9034
rect 7644 8736 8044 8798
rect 7644 8672 7652 8736
rect 7716 8672 7732 8736
rect 7796 8672 7812 8736
rect 7876 8672 7892 8736
rect 7956 8672 7972 8736
rect 8036 8672 8044 8736
rect 7644 7648 8044 8672
rect 7644 7584 7652 7648
rect 7716 7584 7732 7648
rect 7796 7584 7812 7648
rect 7876 7584 7892 7648
rect 7956 7584 7972 7648
rect 8036 7584 8044 7648
rect 7644 6560 8044 7584
rect 7644 6496 7652 6560
rect 7716 6496 7732 6560
rect 7796 6496 7812 6560
rect 7876 6496 7892 6560
rect 7956 6496 7972 6560
rect 8036 6496 8044 6560
rect 7644 5472 8044 6496
rect 7644 5408 7652 5472
rect 7716 5408 7732 5472
rect 7796 5408 7812 5472
rect 7876 5408 7892 5472
rect 7956 5408 7972 5472
rect 8036 5408 8044 5472
rect 7644 5034 8044 5408
rect 7644 4798 7726 5034
rect 7962 4798 8044 5034
rect 7644 4384 8044 4798
rect 7644 4320 7652 4384
rect 7716 4320 7732 4384
rect 7796 4320 7812 4384
rect 7876 4320 7892 4384
rect 7956 4320 7972 4384
rect 8036 4320 8044 4384
rect 7644 3296 8044 4320
rect 7644 3232 7652 3296
rect 7716 3232 7732 3296
rect 7796 3232 7812 3296
rect 7876 3232 7892 3296
rect 7956 3232 7972 3296
rect 8036 3232 8044 3296
rect 7644 2208 8044 3232
rect 7644 2144 7652 2208
rect 7716 2144 7732 2208
rect 7796 2144 7812 2208
rect 7876 2144 7892 2208
rect 7956 2144 7972 2208
rect 8036 2144 8044 2208
rect 7644 2128 8044 2144
rect 10904 10368 11304 11392
rect 10904 10304 10912 10368
rect 10976 10304 10992 10368
rect 11056 10304 11072 10368
rect 11136 10304 11152 10368
rect 11216 10304 11232 10368
rect 11296 10304 11304 10368
rect 10904 9280 11304 10304
rect 10904 9216 10912 9280
rect 10976 9216 10992 9280
rect 11056 9216 11072 9280
rect 11136 9216 11152 9280
rect 11216 9216 11232 9280
rect 11296 9216 11304 9280
rect 10904 8294 11304 9216
rect 10904 8192 10986 8294
rect 11222 8192 11304 8294
rect 10904 8128 10912 8192
rect 10976 8128 10986 8192
rect 11222 8128 11232 8192
rect 11296 8128 11304 8192
rect 10904 8058 10986 8128
rect 11222 8058 11304 8128
rect 10904 7104 11304 8058
rect 10904 7040 10912 7104
rect 10976 7040 10992 7104
rect 11056 7040 11072 7104
rect 11136 7040 11152 7104
rect 11216 7040 11232 7104
rect 11296 7040 11304 7104
rect 10904 6016 11304 7040
rect 10904 5952 10912 6016
rect 10976 5952 10992 6016
rect 11056 5952 11072 6016
rect 11136 5952 11152 6016
rect 11216 5952 11232 6016
rect 11296 5952 11304 6016
rect 10904 4928 11304 5952
rect 10904 4864 10912 4928
rect 10976 4864 10992 4928
rect 11056 4864 11072 4928
rect 11136 4864 11152 4928
rect 11216 4864 11232 4928
rect 11296 4864 11304 4928
rect 10904 4294 11304 4864
rect 10904 4058 10986 4294
rect 11222 4058 11304 4294
rect 10904 3840 11304 4058
rect 10904 3776 10912 3840
rect 10976 3776 10992 3840
rect 11056 3776 11072 3840
rect 11136 3776 11152 3840
rect 11216 3776 11232 3840
rect 11296 3776 11304 3840
rect 10904 2752 11304 3776
rect 10904 2688 10912 2752
rect 10976 2688 10992 2752
rect 11056 2688 11072 2752
rect 11136 2688 11152 2752
rect 11216 2688 11232 2752
rect 11296 2688 11304 2752
rect 10904 2128 11304 2688
rect 11644 27232 12044 27792
rect 11644 27168 11652 27232
rect 11716 27168 11732 27232
rect 11796 27168 11812 27232
rect 11876 27168 11892 27232
rect 11956 27168 11972 27232
rect 12036 27168 12044 27232
rect 11644 26144 12044 27168
rect 11644 26080 11652 26144
rect 11716 26080 11732 26144
rect 11796 26080 11812 26144
rect 11876 26080 11892 26144
rect 11956 26080 11972 26144
rect 12036 26080 12044 26144
rect 11644 25056 12044 26080
rect 11644 24992 11652 25056
rect 11716 25034 11732 25056
rect 11796 25034 11812 25056
rect 11876 25034 11892 25056
rect 11956 25034 11972 25056
rect 11716 24992 11726 25034
rect 11962 24992 11972 25034
rect 12036 24992 12044 25056
rect 11644 24798 11726 24992
rect 11962 24798 12044 24992
rect 11644 23968 12044 24798
rect 11644 23904 11652 23968
rect 11716 23904 11732 23968
rect 11796 23904 11812 23968
rect 11876 23904 11892 23968
rect 11956 23904 11972 23968
rect 12036 23904 12044 23968
rect 11644 22880 12044 23904
rect 11644 22816 11652 22880
rect 11716 22816 11732 22880
rect 11796 22816 11812 22880
rect 11876 22816 11892 22880
rect 11956 22816 11972 22880
rect 12036 22816 12044 22880
rect 11644 21792 12044 22816
rect 11644 21728 11652 21792
rect 11716 21728 11732 21792
rect 11796 21728 11812 21792
rect 11876 21728 11892 21792
rect 11956 21728 11972 21792
rect 12036 21728 12044 21792
rect 11644 21034 12044 21728
rect 11644 20798 11726 21034
rect 11962 20798 12044 21034
rect 11644 20704 12044 20798
rect 11644 20640 11652 20704
rect 11716 20640 11732 20704
rect 11796 20640 11812 20704
rect 11876 20640 11892 20704
rect 11956 20640 11972 20704
rect 12036 20640 12044 20704
rect 11644 19616 12044 20640
rect 11644 19552 11652 19616
rect 11716 19552 11732 19616
rect 11796 19552 11812 19616
rect 11876 19552 11892 19616
rect 11956 19552 11972 19616
rect 12036 19552 12044 19616
rect 11644 18528 12044 19552
rect 11644 18464 11652 18528
rect 11716 18464 11732 18528
rect 11796 18464 11812 18528
rect 11876 18464 11892 18528
rect 11956 18464 11972 18528
rect 12036 18464 12044 18528
rect 11644 17440 12044 18464
rect 14904 27776 15304 27792
rect 14904 27712 14912 27776
rect 14976 27712 14992 27776
rect 15056 27712 15072 27776
rect 15136 27712 15152 27776
rect 15216 27712 15232 27776
rect 15296 27712 15304 27776
rect 14904 26688 15304 27712
rect 14904 26624 14912 26688
rect 14976 26624 14992 26688
rect 15056 26624 15072 26688
rect 15136 26624 15152 26688
rect 15216 26624 15232 26688
rect 15296 26624 15304 26688
rect 14904 25600 15304 26624
rect 14904 25536 14912 25600
rect 14976 25536 14992 25600
rect 15056 25536 15072 25600
rect 15136 25536 15152 25600
rect 15216 25536 15232 25600
rect 15296 25536 15304 25600
rect 14904 24512 15304 25536
rect 14904 24448 14912 24512
rect 14976 24448 14992 24512
rect 15056 24448 15072 24512
rect 15136 24448 15152 24512
rect 15216 24448 15232 24512
rect 15296 24448 15304 24512
rect 14904 24294 15304 24448
rect 14904 24058 14986 24294
rect 15222 24058 15304 24294
rect 14904 23424 15304 24058
rect 14904 23360 14912 23424
rect 14976 23360 14992 23424
rect 15056 23360 15072 23424
rect 15136 23360 15152 23424
rect 15216 23360 15232 23424
rect 15296 23360 15304 23424
rect 14904 22336 15304 23360
rect 14904 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15072 22336
rect 15136 22272 15152 22336
rect 15216 22272 15232 22336
rect 15296 22272 15304 22336
rect 14904 21248 15304 22272
rect 14904 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15072 21248
rect 15136 21184 15152 21248
rect 15216 21184 15232 21248
rect 15296 21184 15304 21248
rect 14904 20294 15304 21184
rect 14904 20160 14986 20294
rect 15222 20160 15304 20294
rect 14904 20096 14912 20160
rect 14976 20096 14986 20160
rect 15222 20096 15232 20160
rect 15296 20096 15304 20160
rect 14904 20058 14986 20096
rect 15222 20058 15304 20096
rect 14904 19072 15304 20058
rect 14904 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15072 19072
rect 15136 19008 15152 19072
rect 15216 19008 15232 19072
rect 15296 19008 15304 19072
rect 14595 18188 14661 18189
rect 14595 18124 14596 18188
rect 14660 18124 14661 18188
rect 14595 18123 14661 18124
rect 11644 17376 11652 17440
rect 11716 17376 11732 17440
rect 11796 17376 11812 17440
rect 11876 17376 11892 17440
rect 11956 17376 11972 17440
rect 12036 17376 12044 17440
rect 11644 17034 12044 17376
rect 11644 16798 11726 17034
rect 11962 16798 12044 17034
rect 11644 16352 12044 16798
rect 11644 16288 11652 16352
rect 11716 16288 11732 16352
rect 11796 16288 11812 16352
rect 11876 16288 11892 16352
rect 11956 16288 11972 16352
rect 12036 16288 12044 16352
rect 11644 15264 12044 16288
rect 14598 16149 14658 18123
rect 14904 17984 15304 19008
rect 14904 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15072 17984
rect 15136 17920 15152 17984
rect 15216 17920 15232 17984
rect 15296 17920 15304 17984
rect 14904 16896 15304 17920
rect 14904 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15072 16896
rect 15136 16832 15152 16896
rect 15216 16832 15232 16896
rect 15296 16832 15304 16896
rect 14904 16294 15304 16832
rect 15644 27232 16044 27792
rect 15644 27168 15652 27232
rect 15716 27168 15732 27232
rect 15796 27168 15812 27232
rect 15876 27168 15892 27232
rect 15956 27168 15972 27232
rect 16036 27168 16044 27232
rect 15644 26144 16044 27168
rect 15644 26080 15652 26144
rect 15716 26080 15732 26144
rect 15796 26080 15812 26144
rect 15876 26080 15892 26144
rect 15956 26080 15972 26144
rect 16036 26080 16044 26144
rect 15644 25056 16044 26080
rect 15644 24992 15652 25056
rect 15716 25034 15732 25056
rect 15796 25034 15812 25056
rect 15876 25034 15892 25056
rect 15956 25034 15972 25056
rect 15716 24992 15726 25034
rect 15962 24992 15972 25034
rect 16036 24992 16044 25056
rect 15644 24798 15726 24992
rect 15962 24798 16044 24992
rect 18904 27776 19304 27792
rect 18904 27712 18912 27776
rect 18976 27712 18992 27776
rect 19056 27712 19072 27776
rect 19136 27712 19152 27776
rect 19216 27712 19232 27776
rect 19296 27712 19304 27776
rect 18904 26688 19304 27712
rect 18904 26624 18912 26688
rect 18976 26624 18992 26688
rect 19056 26624 19072 26688
rect 19136 26624 19152 26688
rect 19216 26624 19232 26688
rect 19296 26624 19304 26688
rect 18904 25600 19304 26624
rect 18904 25536 18912 25600
rect 18976 25536 18992 25600
rect 19056 25536 19072 25600
rect 19136 25536 19152 25600
rect 19216 25536 19232 25600
rect 19296 25536 19304 25600
rect 17539 24988 17605 24989
rect 17539 24924 17540 24988
rect 17604 24924 17605 24988
rect 17539 24923 17605 24924
rect 15644 23968 16044 24798
rect 15644 23904 15652 23968
rect 15716 23904 15732 23968
rect 15796 23904 15812 23968
rect 15876 23904 15892 23968
rect 15956 23904 15972 23968
rect 16036 23904 16044 23968
rect 15644 22880 16044 23904
rect 15644 22816 15652 22880
rect 15716 22816 15732 22880
rect 15796 22816 15812 22880
rect 15876 22816 15892 22880
rect 15956 22816 15972 22880
rect 16036 22816 16044 22880
rect 15644 21792 16044 22816
rect 17355 22540 17421 22541
rect 17355 22476 17356 22540
rect 17420 22476 17421 22540
rect 17355 22475 17421 22476
rect 15644 21728 15652 21792
rect 15716 21728 15732 21792
rect 15796 21728 15812 21792
rect 15876 21728 15892 21792
rect 15956 21728 15972 21792
rect 16036 21728 16044 21792
rect 15644 21034 16044 21728
rect 15644 20798 15726 21034
rect 15962 20798 16044 21034
rect 15644 20704 16044 20798
rect 15644 20640 15652 20704
rect 15716 20640 15732 20704
rect 15796 20640 15812 20704
rect 15876 20640 15892 20704
rect 15956 20640 15972 20704
rect 16036 20640 16044 20704
rect 15644 19616 16044 20640
rect 15644 19552 15652 19616
rect 15716 19552 15732 19616
rect 15796 19552 15812 19616
rect 15876 19552 15892 19616
rect 15956 19552 15972 19616
rect 16036 19552 16044 19616
rect 15644 18528 16044 19552
rect 15644 18464 15652 18528
rect 15716 18464 15732 18528
rect 15796 18464 15812 18528
rect 15876 18464 15892 18528
rect 15956 18464 15972 18528
rect 16036 18464 16044 18528
rect 15644 17440 16044 18464
rect 15644 17376 15652 17440
rect 15716 17376 15732 17440
rect 15796 17376 15812 17440
rect 15876 17376 15892 17440
rect 15956 17376 15972 17440
rect 16036 17376 16044 17440
rect 15644 17034 16044 17376
rect 15644 16798 15726 17034
rect 15962 16798 16044 17034
rect 15515 16692 15581 16693
rect 15515 16628 15516 16692
rect 15580 16628 15581 16692
rect 15515 16627 15581 16628
rect 14595 16148 14661 16149
rect 14595 16084 14596 16148
rect 14660 16084 14661 16148
rect 14595 16083 14661 16084
rect 11644 15200 11652 15264
rect 11716 15200 11732 15264
rect 11796 15200 11812 15264
rect 11876 15200 11892 15264
rect 11956 15200 11972 15264
rect 12036 15200 12044 15264
rect 11644 14176 12044 15200
rect 14598 14517 14658 16083
rect 14904 16058 14986 16294
rect 15222 16058 15304 16294
rect 14904 15808 15304 16058
rect 14904 15744 14912 15808
rect 14976 15744 14992 15808
rect 15056 15744 15072 15808
rect 15136 15744 15152 15808
rect 15216 15744 15232 15808
rect 15296 15744 15304 15808
rect 14904 14720 15304 15744
rect 14904 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15072 14720
rect 15136 14656 15152 14720
rect 15216 14656 15232 14720
rect 15296 14656 15304 14720
rect 14595 14516 14661 14517
rect 14595 14452 14596 14516
rect 14660 14452 14661 14516
rect 14595 14451 14661 14452
rect 11644 14112 11652 14176
rect 11716 14112 11732 14176
rect 11796 14112 11812 14176
rect 11876 14112 11892 14176
rect 11956 14112 11972 14176
rect 12036 14112 12044 14176
rect 11644 13088 12044 14112
rect 11644 13024 11652 13088
rect 11716 13034 11732 13088
rect 11796 13034 11812 13088
rect 11876 13034 11892 13088
rect 11956 13034 11972 13088
rect 11716 13024 11726 13034
rect 11962 13024 11972 13034
rect 12036 13024 12044 13088
rect 11644 12798 11726 13024
rect 11962 12798 12044 13024
rect 11644 12000 12044 12798
rect 11644 11936 11652 12000
rect 11716 11936 11732 12000
rect 11796 11936 11812 12000
rect 11876 11936 11892 12000
rect 11956 11936 11972 12000
rect 12036 11936 12044 12000
rect 11644 10912 12044 11936
rect 11644 10848 11652 10912
rect 11716 10848 11732 10912
rect 11796 10848 11812 10912
rect 11876 10848 11892 10912
rect 11956 10848 11972 10912
rect 12036 10848 12044 10912
rect 11644 9824 12044 10848
rect 11644 9760 11652 9824
rect 11716 9760 11732 9824
rect 11796 9760 11812 9824
rect 11876 9760 11892 9824
rect 11956 9760 11972 9824
rect 12036 9760 12044 9824
rect 11644 9034 12044 9760
rect 11644 8798 11726 9034
rect 11962 8798 12044 9034
rect 11644 8736 12044 8798
rect 11644 8672 11652 8736
rect 11716 8672 11732 8736
rect 11796 8672 11812 8736
rect 11876 8672 11892 8736
rect 11956 8672 11972 8736
rect 12036 8672 12044 8736
rect 11644 7648 12044 8672
rect 14598 8533 14658 14451
rect 14904 13632 15304 14656
rect 15518 14517 15578 16627
rect 15644 16352 16044 16798
rect 15644 16288 15652 16352
rect 15716 16288 15732 16352
rect 15796 16288 15812 16352
rect 15876 16288 15892 16352
rect 15956 16288 15972 16352
rect 16036 16288 16044 16352
rect 15644 15264 16044 16288
rect 15644 15200 15652 15264
rect 15716 15200 15732 15264
rect 15796 15200 15812 15264
rect 15876 15200 15892 15264
rect 15956 15200 15972 15264
rect 16036 15200 16044 15264
rect 15515 14516 15581 14517
rect 15515 14452 15516 14516
rect 15580 14452 15581 14516
rect 15515 14451 15581 14452
rect 14904 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15072 13632
rect 15136 13568 15152 13632
rect 15216 13568 15232 13632
rect 15296 13568 15304 13632
rect 14904 12544 15304 13568
rect 14904 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15072 12544
rect 15136 12480 15152 12544
rect 15216 12480 15232 12544
rect 15296 12480 15304 12544
rect 14904 12294 15304 12480
rect 14904 12058 14986 12294
rect 15222 12058 15304 12294
rect 14904 11456 15304 12058
rect 14904 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15072 11456
rect 15136 11392 15152 11456
rect 15216 11392 15232 11456
rect 15296 11392 15304 11456
rect 14904 10368 15304 11392
rect 14904 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15072 10368
rect 15136 10304 15152 10368
rect 15216 10304 15232 10368
rect 15296 10304 15304 10368
rect 14904 9280 15304 10304
rect 14904 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15072 9280
rect 15136 9216 15152 9280
rect 15216 9216 15232 9280
rect 15296 9216 15304 9280
rect 14595 8532 14661 8533
rect 14595 8468 14596 8532
rect 14660 8468 14661 8532
rect 14595 8467 14661 8468
rect 11644 7584 11652 7648
rect 11716 7584 11732 7648
rect 11796 7584 11812 7648
rect 11876 7584 11892 7648
rect 11956 7584 11972 7648
rect 12036 7584 12044 7648
rect 11644 6560 12044 7584
rect 11644 6496 11652 6560
rect 11716 6496 11732 6560
rect 11796 6496 11812 6560
rect 11876 6496 11892 6560
rect 11956 6496 11972 6560
rect 12036 6496 12044 6560
rect 11644 5472 12044 6496
rect 11644 5408 11652 5472
rect 11716 5408 11732 5472
rect 11796 5408 11812 5472
rect 11876 5408 11892 5472
rect 11956 5408 11972 5472
rect 12036 5408 12044 5472
rect 11644 5034 12044 5408
rect 11644 4798 11726 5034
rect 11962 4798 12044 5034
rect 11644 4384 12044 4798
rect 11644 4320 11652 4384
rect 11716 4320 11732 4384
rect 11796 4320 11812 4384
rect 11876 4320 11892 4384
rect 11956 4320 11972 4384
rect 12036 4320 12044 4384
rect 11644 3296 12044 4320
rect 11644 3232 11652 3296
rect 11716 3232 11732 3296
rect 11796 3232 11812 3296
rect 11876 3232 11892 3296
rect 11956 3232 11972 3296
rect 12036 3232 12044 3296
rect 11644 2208 12044 3232
rect 11644 2144 11652 2208
rect 11716 2144 11732 2208
rect 11796 2144 11812 2208
rect 11876 2144 11892 2208
rect 11956 2144 11972 2208
rect 12036 2144 12044 2208
rect 11644 2128 12044 2144
rect 14904 8294 15304 9216
rect 14904 8192 14986 8294
rect 15222 8192 15304 8294
rect 14904 8128 14912 8192
rect 14976 8128 14986 8192
rect 15222 8128 15232 8192
rect 15296 8128 15304 8192
rect 14904 8058 14986 8128
rect 15222 8058 15304 8128
rect 14904 7104 15304 8058
rect 14904 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15072 7104
rect 15136 7040 15152 7104
rect 15216 7040 15232 7104
rect 15296 7040 15304 7104
rect 14904 6016 15304 7040
rect 14904 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15072 6016
rect 15136 5952 15152 6016
rect 15216 5952 15232 6016
rect 15296 5952 15304 6016
rect 14904 4928 15304 5952
rect 14904 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15072 4928
rect 15136 4864 15152 4928
rect 15216 4864 15232 4928
rect 15296 4864 15304 4928
rect 14904 4294 15304 4864
rect 14904 4058 14986 4294
rect 15222 4058 15304 4294
rect 14904 3840 15304 4058
rect 14904 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15072 3840
rect 15136 3776 15152 3840
rect 15216 3776 15232 3840
rect 15296 3776 15304 3840
rect 14904 2752 15304 3776
rect 14904 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15072 2752
rect 15136 2688 15152 2752
rect 15216 2688 15232 2752
rect 15296 2688 15304 2752
rect 14904 2128 15304 2688
rect 15644 14176 16044 15200
rect 15644 14112 15652 14176
rect 15716 14112 15732 14176
rect 15796 14112 15812 14176
rect 15876 14112 15892 14176
rect 15956 14112 15972 14176
rect 16036 14112 16044 14176
rect 15644 13088 16044 14112
rect 15644 13024 15652 13088
rect 15716 13034 15732 13088
rect 15796 13034 15812 13088
rect 15876 13034 15892 13088
rect 15956 13034 15972 13088
rect 15716 13024 15726 13034
rect 15962 13024 15972 13034
rect 16036 13024 16044 13088
rect 15644 12798 15726 13024
rect 15962 12798 16044 13024
rect 15644 12000 16044 12798
rect 15644 11936 15652 12000
rect 15716 11936 15732 12000
rect 15796 11936 15812 12000
rect 15876 11936 15892 12000
rect 15956 11936 15972 12000
rect 16036 11936 16044 12000
rect 15644 10912 16044 11936
rect 15644 10848 15652 10912
rect 15716 10848 15732 10912
rect 15796 10848 15812 10912
rect 15876 10848 15892 10912
rect 15956 10848 15972 10912
rect 16036 10848 16044 10912
rect 15644 9824 16044 10848
rect 17358 10709 17418 22475
rect 17355 10708 17421 10709
rect 17355 10644 17356 10708
rect 17420 10644 17421 10708
rect 17355 10643 17421 10644
rect 17542 10301 17602 24923
rect 18904 24512 19304 25536
rect 18904 24448 18912 24512
rect 18976 24448 18992 24512
rect 19056 24448 19072 24512
rect 19136 24448 19152 24512
rect 19216 24448 19232 24512
rect 19296 24448 19304 24512
rect 18904 24294 19304 24448
rect 18904 24058 18986 24294
rect 19222 24058 19304 24294
rect 18904 23424 19304 24058
rect 18904 23360 18912 23424
rect 18976 23360 18992 23424
rect 19056 23360 19072 23424
rect 19136 23360 19152 23424
rect 19216 23360 19232 23424
rect 19296 23360 19304 23424
rect 18904 22336 19304 23360
rect 18904 22272 18912 22336
rect 18976 22272 18992 22336
rect 19056 22272 19072 22336
rect 19136 22272 19152 22336
rect 19216 22272 19232 22336
rect 19296 22272 19304 22336
rect 18904 21248 19304 22272
rect 18904 21184 18912 21248
rect 18976 21184 18992 21248
rect 19056 21184 19072 21248
rect 19136 21184 19152 21248
rect 19216 21184 19232 21248
rect 19296 21184 19304 21248
rect 18275 20364 18341 20365
rect 18275 20300 18276 20364
rect 18340 20300 18341 20364
rect 18275 20299 18341 20300
rect 18278 14381 18338 20299
rect 18904 20294 19304 21184
rect 19644 27232 20044 27792
rect 19644 27168 19652 27232
rect 19716 27168 19732 27232
rect 19796 27168 19812 27232
rect 19876 27168 19892 27232
rect 19956 27168 19972 27232
rect 20036 27168 20044 27232
rect 19644 26144 20044 27168
rect 19644 26080 19652 26144
rect 19716 26080 19732 26144
rect 19796 26080 19812 26144
rect 19876 26080 19892 26144
rect 19956 26080 19972 26144
rect 20036 26080 20044 26144
rect 19644 25056 20044 26080
rect 19644 24992 19652 25056
rect 19716 25034 19732 25056
rect 19796 25034 19812 25056
rect 19876 25034 19892 25056
rect 19956 25034 19972 25056
rect 19716 24992 19726 25034
rect 19962 24992 19972 25034
rect 20036 24992 20044 25056
rect 19644 24798 19726 24992
rect 19962 24798 20044 24992
rect 19644 23968 20044 24798
rect 19644 23904 19652 23968
rect 19716 23904 19732 23968
rect 19796 23904 19812 23968
rect 19876 23904 19892 23968
rect 19956 23904 19972 23968
rect 20036 23904 20044 23968
rect 19644 22880 20044 23904
rect 19644 22816 19652 22880
rect 19716 22816 19732 22880
rect 19796 22816 19812 22880
rect 19876 22816 19892 22880
rect 19956 22816 19972 22880
rect 20036 22816 20044 22880
rect 19644 21792 20044 22816
rect 19644 21728 19652 21792
rect 19716 21728 19732 21792
rect 19796 21728 19812 21792
rect 19876 21728 19892 21792
rect 19956 21728 19972 21792
rect 20036 21728 20044 21792
rect 19644 21034 20044 21728
rect 19379 20908 19445 20909
rect 19379 20844 19380 20908
rect 19444 20844 19445 20908
rect 19379 20843 19445 20844
rect 18904 20160 18986 20294
rect 19222 20160 19304 20294
rect 18904 20096 18912 20160
rect 18976 20096 18986 20160
rect 19222 20096 19232 20160
rect 19296 20096 19304 20160
rect 18904 20058 18986 20096
rect 19222 20058 19304 20096
rect 18904 19072 19304 20058
rect 18904 19008 18912 19072
rect 18976 19008 18992 19072
rect 19056 19008 19072 19072
rect 19136 19008 19152 19072
rect 19216 19008 19232 19072
rect 19296 19008 19304 19072
rect 18904 17984 19304 19008
rect 18904 17920 18912 17984
rect 18976 17920 18992 17984
rect 19056 17920 19072 17984
rect 19136 17920 19152 17984
rect 19216 17920 19232 17984
rect 19296 17920 19304 17984
rect 18904 16896 19304 17920
rect 18904 16832 18912 16896
rect 18976 16832 18992 16896
rect 19056 16832 19072 16896
rect 19136 16832 19152 16896
rect 19216 16832 19232 16896
rect 19296 16832 19304 16896
rect 18904 16294 19304 16832
rect 18643 16284 18709 16285
rect 18643 16220 18644 16284
rect 18708 16220 18709 16284
rect 18643 16219 18709 16220
rect 18275 14380 18341 14381
rect 18275 14316 18276 14380
rect 18340 14316 18341 14380
rect 18275 14315 18341 14316
rect 18278 10301 18338 14315
rect 18459 13428 18525 13429
rect 18459 13364 18460 13428
rect 18524 13364 18525 13428
rect 18459 13363 18525 13364
rect 17539 10300 17605 10301
rect 17539 10236 17540 10300
rect 17604 10236 17605 10300
rect 17539 10235 17605 10236
rect 18275 10300 18341 10301
rect 18275 10236 18276 10300
rect 18340 10236 18341 10300
rect 18275 10235 18341 10236
rect 15644 9760 15652 9824
rect 15716 9760 15732 9824
rect 15796 9760 15812 9824
rect 15876 9760 15892 9824
rect 15956 9760 15972 9824
rect 16036 9760 16044 9824
rect 15644 9034 16044 9760
rect 15644 8798 15726 9034
rect 15962 8798 16044 9034
rect 15644 8736 16044 8798
rect 15644 8672 15652 8736
rect 15716 8672 15732 8736
rect 15796 8672 15812 8736
rect 15876 8672 15892 8736
rect 15956 8672 15972 8736
rect 16036 8672 16044 8736
rect 15644 7648 16044 8672
rect 15644 7584 15652 7648
rect 15716 7584 15732 7648
rect 15796 7584 15812 7648
rect 15876 7584 15892 7648
rect 15956 7584 15972 7648
rect 16036 7584 16044 7648
rect 15644 6560 16044 7584
rect 18462 6765 18522 13363
rect 18646 7989 18706 16219
rect 18904 16058 18986 16294
rect 19222 16058 19304 16294
rect 19382 16285 19442 20843
rect 19644 20798 19726 21034
rect 19962 20798 20044 21034
rect 19644 20704 20044 20798
rect 19644 20640 19652 20704
rect 19716 20640 19732 20704
rect 19796 20640 19812 20704
rect 19876 20640 19892 20704
rect 19956 20640 19972 20704
rect 20036 20640 20044 20704
rect 19644 19616 20044 20640
rect 19644 19552 19652 19616
rect 19716 19552 19732 19616
rect 19796 19552 19812 19616
rect 19876 19552 19892 19616
rect 19956 19552 19972 19616
rect 20036 19552 20044 19616
rect 19644 18528 20044 19552
rect 19644 18464 19652 18528
rect 19716 18464 19732 18528
rect 19796 18464 19812 18528
rect 19876 18464 19892 18528
rect 19956 18464 19972 18528
rect 20036 18464 20044 18528
rect 19644 17440 20044 18464
rect 19644 17376 19652 17440
rect 19716 17376 19732 17440
rect 19796 17376 19812 17440
rect 19876 17376 19892 17440
rect 19956 17376 19972 17440
rect 20036 17376 20044 17440
rect 19644 17034 20044 17376
rect 19644 16798 19726 17034
rect 19962 16798 20044 17034
rect 19644 16352 20044 16798
rect 19644 16288 19652 16352
rect 19716 16288 19732 16352
rect 19796 16288 19812 16352
rect 19876 16288 19892 16352
rect 19956 16288 19972 16352
rect 20036 16288 20044 16352
rect 19379 16284 19445 16285
rect 19379 16220 19380 16284
rect 19444 16220 19445 16284
rect 19379 16219 19445 16220
rect 18904 15808 19304 16058
rect 18904 15744 18912 15808
rect 18976 15744 18992 15808
rect 19056 15744 19072 15808
rect 19136 15744 19152 15808
rect 19216 15744 19232 15808
rect 19296 15744 19304 15808
rect 18904 14720 19304 15744
rect 18904 14656 18912 14720
rect 18976 14656 18992 14720
rect 19056 14656 19072 14720
rect 19136 14656 19152 14720
rect 19216 14656 19232 14720
rect 19296 14656 19304 14720
rect 18904 13632 19304 14656
rect 18904 13568 18912 13632
rect 18976 13568 18992 13632
rect 19056 13568 19072 13632
rect 19136 13568 19152 13632
rect 19216 13568 19232 13632
rect 19296 13568 19304 13632
rect 18904 12544 19304 13568
rect 18904 12480 18912 12544
rect 18976 12480 18992 12544
rect 19056 12480 19072 12544
rect 19136 12480 19152 12544
rect 19216 12480 19232 12544
rect 19296 12480 19304 12544
rect 18904 12294 19304 12480
rect 18904 12058 18986 12294
rect 19222 12058 19304 12294
rect 18904 11456 19304 12058
rect 18904 11392 18912 11456
rect 18976 11392 18992 11456
rect 19056 11392 19072 11456
rect 19136 11392 19152 11456
rect 19216 11392 19232 11456
rect 19296 11392 19304 11456
rect 18904 10368 19304 11392
rect 18904 10304 18912 10368
rect 18976 10304 18992 10368
rect 19056 10304 19072 10368
rect 19136 10304 19152 10368
rect 19216 10304 19232 10368
rect 19296 10304 19304 10368
rect 18904 9280 19304 10304
rect 18904 9216 18912 9280
rect 18976 9216 18992 9280
rect 19056 9216 19072 9280
rect 19136 9216 19152 9280
rect 19216 9216 19232 9280
rect 19296 9216 19304 9280
rect 18904 8294 19304 9216
rect 18904 8192 18986 8294
rect 19222 8192 19304 8294
rect 18904 8128 18912 8192
rect 18976 8128 18986 8192
rect 19222 8128 19232 8192
rect 19296 8128 19304 8192
rect 18904 8058 18986 8128
rect 19222 8058 19304 8128
rect 18643 7988 18709 7989
rect 18643 7924 18644 7988
rect 18708 7924 18709 7988
rect 18643 7923 18709 7924
rect 18904 7104 19304 8058
rect 18904 7040 18912 7104
rect 18976 7040 18992 7104
rect 19056 7040 19072 7104
rect 19136 7040 19152 7104
rect 19216 7040 19232 7104
rect 19296 7040 19304 7104
rect 18459 6764 18525 6765
rect 18459 6700 18460 6764
rect 18524 6700 18525 6764
rect 18459 6699 18525 6700
rect 15644 6496 15652 6560
rect 15716 6496 15732 6560
rect 15796 6496 15812 6560
rect 15876 6496 15892 6560
rect 15956 6496 15972 6560
rect 16036 6496 16044 6560
rect 15644 5472 16044 6496
rect 15644 5408 15652 5472
rect 15716 5408 15732 5472
rect 15796 5408 15812 5472
rect 15876 5408 15892 5472
rect 15956 5408 15972 5472
rect 16036 5408 16044 5472
rect 15644 5034 16044 5408
rect 15644 4798 15726 5034
rect 15962 4798 16044 5034
rect 15644 4384 16044 4798
rect 15644 4320 15652 4384
rect 15716 4320 15732 4384
rect 15796 4320 15812 4384
rect 15876 4320 15892 4384
rect 15956 4320 15972 4384
rect 16036 4320 16044 4384
rect 15644 3296 16044 4320
rect 15644 3232 15652 3296
rect 15716 3232 15732 3296
rect 15796 3232 15812 3296
rect 15876 3232 15892 3296
rect 15956 3232 15972 3296
rect 16036 3232 16044 3296
rect 15644 2208 16044 3232
rect 15644 2144 15652 2208
rect 15716 2144 15732 2208
rect 15796 2144 15812 2208
rect 15876 2144 15892 2208
rect 15956 2144 15972 2208
rect 16036 2144 16044 2208
rect 15644 2128 16044 2144
rect 18904 6016 19304 7040
rect 18904 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19304 6016
rect 18904 4928 19304 5952
rect 18904 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19304 4928
rect 18904 4294 19304 4864
rect 18904 4058 18986 4294
rect 19222 4058 19304 4294
rect 18904 3840 19304 4058
rect 18904 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19304 3840
rect 18904 2752 19304 3776
rect 18904 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19304 2752
rect 18904 2128 19304 2688
rect 19644 15264 20044 16288
rect 19644 15200 19652 15264
rect 19716 15200 19732 15264
rect 19796 15200 19812 15264
rect 19876 15200 19892 15264
rect 19956 15200 19972 15264
rect 20036 15200 20044 15264
rect 19644 14176 20044 15200
rect 19644 14112 19652 14176
rect 19716 14112 19732 14176
rect 19796 14112 19812 14176
rect 19876 14112 19892 14176
rect 19956 14112 19972 14176
rect 20036 14112 20044 14176
rect 19644 13088 20044 14112
rect 19644 13024 19652 13088
rect 19716 13034 19732 13088
rect 19796 13034 19812 13088
rect 19876 13034 19892 13088
rect 19956 13034 19972 13088
rect 19716 13024 19726 13034
rect 19962 13024 19972 13034
rect 20036 13024 20044 13088
rect 19644 12798 19726 13024
rect 19962 12798 20044 13024
rect 19644 12000 20044 12798
rect 19644 11936 19652 12000
rect 19716 11936 19732 12000
rect 19796 11936 19812 12000
rect 19876 11936 19892 12000
rect 19956 11936 19972 12000
rect 20036 11936 20044 12000
rect 19644 10912 20044 11936
rect 19644 10848 19652 10912
rect 19716 10848 19732 10912
rect 19796 10848 19812 10912
rect 19876 10848 19892 10912
rect 19956 10848 19972 10912
rect 20036 10848 20044 10912
rect 19644 9824 20044 10848
rect 19644 9760 19652 9824
rect 19716 9760 19732 9824
rect 19796 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20044 9824
rect 19644 9034 20044 9760
rect 19644 8798 19726 9034
rect 19962 8798 20044 9034
rect 19644 8736 20044 8798
rect 19644 8672 19652 8736
rect 19716 8672 19732 8736
rect 19796 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20044 8736
rect 19644 7648 20044 8672
rect 19644 7584 19652 7648
rect 19716 7584 19732 7648
rect 19796 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20044 7648
rect 19644 6560 20044 7584
rect 19644 6496 19652 6560
rect 19716 6496 19732 6560
rect 19796 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20044 6560
rect 19644 5472 20044 6496
rect 19644 5408 19652 5472
rect 19716 5408 19732 5472
rect 19796 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20044 5472
rect 19644 5034 20044 5408
rect 19644 4798 19726 5034
rect 19962 4798 20044 5034
rect 19644 4384 20044 4798
rect 19644 4320 19652 4384
rect 19716 4320 19732 4384
rect 19796 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20044 4384
rect 19644 3296 20044 4320
rect 19644 3232 19652 3296
rect 19716 3232 19732 3296
rect 19796 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20044 3296
rect 19644 2208 20044 3232
rect 19644 2144 19652 2208
rect 19716 2144 19732 2208
rect 19796 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20044 2208
rect 19644 2128 20044 2144
rect 22904 27776 23304 27792
rect 22904 27712 22912 27776
rect 22976 27712 22992 27776
rect 23056 27712 23072 27776
rect 23136 27712 23152 27776
rect 23216 27712 23232 27776
rect 23296 27712 23304 27776
rect 22904 26688 23304 27712
rect 22904 26624 22912 26688
rect 22976 26624 22992 26688
rect 23056 26624 23072 26688
rect 23136 26624 23152 26688
rect 23216 26624 23232 26688
rect 23296 26624 23304 26688
rect 22904 25600 23304 26624
rect 22904 25536 22912 25600
rect 22976 25536 22992 25600
rect 23056 25536 23072 25600
rect 23136 25536 23152 25600
rect 23216 25536 23232 25600
rect 23296 25536 23304 25600
rect 22904 24512 23304 25536
rect 22904 24448 22912 24512
rect 22976 24448 22992 24512
rect 23056 24448 23072 24512
rect 23136 24448 23152 24512
rect 23216 24448 23232 24512
rect 23296 24448 23304 24512
rect 22904 24294 23304 24448
rect 22904 24058 22986 24294
rect 23222 24058 23304 24294
rect 22904 23424 23304 24058
rect 22904 23360 22912 23424
rect 22976 23360 22992 23424
rect 23056 23360 23072 23424
rect 23136 23360 23152 23424
rect 23216 23360 23232 23424
rect 23296 23360 23304 23424
rect 22904 22336 23304 23360
rect 22904 22272 22912 22336
rect 22976 22272 22992 22336
rect 23056 22272 23072 22336
rect 23136 22272 23152 22336
rect 23216 22272 23232 22336
rect 23296 22272 23304 22336
rect 22904 21248 23304 22272
rect 22904 21184 22912 21248
rect 22976 21184 22992 21248
rect 23056 21184 23072 21248
rect 23136 21184 23152 21248
rect 23216 21184 23232 21248
rect 23296 21184 23304 21248
rect 22904 20294 23304 21184
rect 22904 20160 22986 20294
rect 23222 20160 23304 20294
rect 22904 20096 22912 20160
rect 22976 20096 22986 20160
rect 23222 20096 23232 20160
rect 23296 20096 23304 20160
rect 22904 20058 22986 20096
rect 23222 20058 23304 20096
rect 22904 19072 23304 20058
rect 22904 19008 22912 19072
rect 22976 19008 22992 19072
rect 23056 19008 23072 19072
rect 23136 19008 23152 19072
rect 23216 19008 23232 19072
rect 23296 19008 23304 19072
rect 22904 17984 23304 19008
rect 22904 17920 22912 17984
rect 22976 17920 22992 17984
rect 23056 17920 23072 17984
rect 23136 17920 23152 17984
rect 23216 17920 23232 17984
rect 23296 17920 23304 17984
rect 22904 16896 23304 17920
rect 22904 16832 22912 16896
rect 22976 16832 22992 16896
rect 23056 16832 23072 16896
rect 23136 16832 23152 16896
rect 23216 16832 23232 16896
rect 23296 16832 23304 16896
rect 22904 16294 23304 16832
rect 22904 16058 22986 16294
rect 23222 16058 23304 16294
rect 22904 15808 23304 16058
rect 22904 15744 22912 15808
rect 22976 15744 22992 15808
rect 23056 15744 23072 15808
rect 23136 15744 23152 15808
rect 23216 15744 23232 15808
rect 23296 15744 23304 15808
rect 22904 14720 23304 15744
rect 22904 14656 22912 14720
rect 22976 14656 22992 14720
rect 23056 14656 23072 14720
rect 23136 14656 23152 14720
rect 23216 14656 23232 14720
rect 23296 14656 23304 14720
rect 22904 13632 23304 14656
rect 22904 13568 22912 13632
rect 22976 13568 22992 13632
rect 23056 13568 23072 13632
rect 23136 13568 23152 13632
rect 23216 13568 23232 13632
rect 23296 13568 23304 13632
rect 22904 12544 23304 13568
rect 22904 12480 22912 12544
rect 22976 12480 22992 12544
rect 23056 12480 23072 12544
rect 23136 12480 23152 12544
rect 23216 12480 23232 12544
rect 23296 12480 23304 12544
rect 22904 12294 23304 12480
rect 22904 12058 22986 12294
rect 23222 12058 23304 12294
rect 22904 11456 23304 12058
rect 22904 11392 22912 11456
rect 22976 11392 22992 11456
rect 23056 11392 23072 11456
rect 23136 11392 23152 11456
rect 23216 11392 23232 11456
rect 23296 11392 23304 11456
rect 22904 10368 23304 11392
rect 22904 10304 22912 10368
rect 22976 10304 22992 10368
rect 23056 10304 23072 10368
rect 23136 10304 23152 10368
rect 23216 10304 23232 10368
rect 23296 10304 23304 10368
rect 22904 9280 23304 10304
rect 22904 9216 22912 9280
rect 22976 9216 22992 9280
rect 23056 9216 23072 9280
rect 23136 9216 23152 9280
rect 23216 9216 23232 9280
rect 23296 9216 23304 9280
rect 22904 8294 23304 9216
rect 22904 8192 22986 8294
rect 23222 8192 23304 8294
rect 22904 8128 22912 8192
rect 22976 8128 22986 8192
rect 23222 8128 23232 8192
rect 23296 8128 23304 8192
rect 22904 8058 22986 8128
rect 23222 8058 23304 8128
rect 22904 7104 23304 8058
rect 22904 7040 22912 7104
rect 22976 7040 22992 7104
rect 23056 7040 23072 7104
rect 23136 7040 23152 7104
rect 23216 7040 23232 7104
rect 23296 7040 23304 7104
rect 22904 6016 23304 7040
rect 22904 5952 22912 6016
rect 22976 5952 22992 6016
rect 23056 5952 23072 6016
rect 23136 5952 23152 6016
rect 23216 5952 23232 6016
rect 23296 5952 23304 6016
rect 22904 4928 23304 5952
rect 22904 4864 22912 4928
rect 22976 4864 22992 4928
rect 23056 4864 23072 4928
rect 23136 4864 23152 4928
rect 23216 4864 23232 4928
rect 23296 4864 23304 4928
rect 22904 4294 23304 4864
rect 22904 4058 22986 4294
rect 23222 4058 23304 4294
rect 22904 3840 23304 4058
rect 22904 3776 22912 3840
rect 22976 3776 22992 3840
rect 23056 3776 23072 3840
rect 23136 3776 23152 3840
rect 23216 3776 23232 3840
rect 23296 3776 23304 3840
rect 22904 2752 23304 3776
rect 22904 2688 22912 2752
rect 22976 2688 22992 2752
rect 23056 2688 23072 2752
rect 23136 2688 23152 2752
rect 23216 2688 23232 2752
rect 23296 2688 23304 2752
rect 22904 2128 23304 2688
rect 23644 27232 24044 27792
rect 23644 27168 23652 27232
rect 23716 27168 23732 27232
rect 23796 27168 23812 27232
rect 23876 27168 23892 27232
rect 23956 27168 23972 27232
rect 24036 27168 24044 27232
rect 23644 26144 24044 27168
rect 23644 26080 23652 26144
rect 23716 26080 23732 26144
rect 23796 26080 23812 26144
rect 23876 26080 23892 26144
rect 23956 26080 23972 26144
rect 24036 26080 24044 26144
rect 23644 25056 24044 26080
rect 23644 24992 23652 25056
rect 23716 25034 23732 25056
rect 23796 25034 23812 25056
rect 23876 25034 23892 25056
rect 23956 25034 23972 25056
rect 23716 24992 23726 25034
rect 23962 24992 23972 25034
rect 24036 24992 24044 25056
rect 23644 24798 23726 24992
rect 23962 24798 24044 24992
rect 24347 24988 24413 24989
rect 24347 24924 24348 24988
rect 24412 24924 24413 24988
rect 24347 24923 24413 24924
rect 23644 23968 24044 24798
rect 23644 23904 23652 23968
rect 23716 23904 23732 23968
rect 23796 23904 23812 23968
rect 23876 23904 23892 23968
rect 23956 23904 23972 23968
rect 24036 23904 24044 23968
rect 23644 22880 24044 23904
rect 23644 22816 23652 22880
rect 23716 22816 23732 22880
rect 23796 22816 23812 22880
rect 23876 22816 23892 22880
rect 23956 22816 23972 22880
rect 24036 22816 24044 22880
rect 23644 21792 24044 22816
rect 24350 21997 24410 24923
rect 24347 21996 24413 21997
rect 24347 21932 24348 21996
rect 24412 21932 24413 21996
rect 24347 21931 24413 21932
rect 23644 21728 23652 21792
rect 23716 21728 23732 21792
rect 23796 21728 23812 21792
rect 23876 21728 23892 21792
rect 23956 21728 23972 21792
rect 24036 21728 24044 21792
rect 23644 21034 24044 21728
rect 23644 20798 23726 21034
rect 23962 20798 24044 21034
rect 23644 20704 24044 20798
rect 23644 20640 23652 20704
rect 23716 20640 23732 20704
rect 23796 20640 23812 20704
rect 23876 20640 23892 20704
rect 23956 20640 23972 20704
rect 24036 20640 24044 20704
rect 23644 19616 24044 20640
rect 23644 19552 23652 19616
rect 23716 19552 23732 19616
rect 23796 19552 23812 19616
rect 23876 19552 23892 19616
rect 23956 19552 23972 19616
rect 24036 19552 24044 19616
rect 23644 18528 24044 19552
rect 23644 18464 23652 18528
rect 23716 18464 23732 18528
rect 23796 18464 23812 18528
rect 23876 18464 23892 18528
rect 23956 18464 23972 18528
rect 24036 18464 24044 18528
rect 23644 17440 24044 18464
rect 23644 17376 23652 17440
rect 23716 17376 23732 17440
rect 23796 17376 23812 17440
rect 23876 17376 23892 17440
rect 23956 17376 23972 17440
rect 24036 17376 24044 17440
rect 23644 17034 24044 17376
rect 23644 16798 23726 17034
rect 23962 16798 24044 17034
rect 23644 16352 24044 16798
rect 23644 16288 23652 16352
rect 23716 16288 23732 16352
rect 23796 16288 23812 16352
rect 23876 16288 23892 16352
rect 23956 16288 23972 16352
rect 24036 16288 24044 16352
rect 23644 15264 24044 16288
rect 23644 15200 23652 15264
rect 23716 15200 23732 15264
rect 23796 15200 23812 15264
rect 23876 15200 23892 15264
rect 23956 15200 23972 15264
rect 24036 15200 24044 15264
rect 23644 14176 24044 15200
rect 23644 14112 23652 14176
rect 23716 14112 23732 14176
rect 23796 14112 23812 14176
rect 23876 14112 23892 14176
rect 23956 14112 23972 14176
rect 24036 14112 24044 14176
rect 23644 13088 24044 14112
rect 23644 13024 23652 13088
rect 23716 13034 23732 13088
rect 23796 13034 23812 13088
rect 23876 13034 23892 13088
rect 23956 13034 23972 13088
rect 23716 13024 23726 13034
rect 23962 13024 23972 13034
rect 24036 13024 24044 13088
rect 23644 12798 23726 13024
rect 23962 12798 24044 13024
rect 23644 12000 24044 12798
rect 23644 11936 23652 12000
rect 23716 11936 23732 12000
rect 23796 11936 23812 12000
rect 23876 11936 23892 12000
rect 23956 11936 23972 12000
rect 24036 11936 24044 12000
rect 23644 10912 24044 11936
rect 23644 10848 23652 10912
rect 23716 10848 23732 10912
rect 23796 10848 23812 10912
rect 23876 10848 23892 10912
rect 23956 10848 23972 10912
rect 24036 10848 24044 10912
rect 23644 9824 24044 10848
rect 23644 9760 23652 9824
rect 23716 9760 23732 9824
rect 23796 9760 23812 9824
rect 23876 9760 23892 9824
rect 23956 9760 23972 9824
rect 24036 9760 24044 9824
rect 23644 9034 24044 9760
rect 23644 8798 23726 9034
rect 23962 8798 24044 9034
rect 23644 8736 24044 8798
rect 23644 8672 23652 8736
rect 23716 8672 23732 8736
rect 23796 8672 23812 8736
rect 23876 8672 23892 8736
rect 23956 8672 23972 8736
rect 24036 8672 24044 8736
rect 23644 7648 24044 8672
rect 23644 7584 23652 7648
rect 23716 7584 23732 7648
rect 23796 7584 23812 7648
rect 23876 7584 23892 7648
rect 23956 7584 23972 7648
rect 24036 7584 24044 7648
rect 23644 6560 24044 7584
rect 23644 6496 23652 6560
rect 23716 6496 23732 6560
rect 23796 6496 23812 6560
rect 23876 6496 23892 6560
rect 23956 6496 23972 6560
rect 24036 6496 24044 6560
rect 23644 5472 24044 6496
rect 23644 5408 23652 5472
rect 23716 5408 23732 5472
rect 23796 5408 23812 5472
rect 23876 5408 23892 5472
rect 23956 5408 23972 5472
rect 24036 5408 24044 5472
rect 23644 5034 24044 5408
rect 23644 4798 23726 5034
rect 23962 4798 24044 5034
rect 23644 4384 24044 4798
rect 23644 4320 23652 4384
rect 23716 4320 23732 4384
rect 23796 4320 23812 4384
rect 23876 4320 23892 4384
rect 23956 4320 23972 4384
rect 24036 4320 24044 4384
rect 23644 3296 24044 4320
rect 23644 3232 23652 3296
rect 23716 3232 23732 3296
rect 23796 3232 23812 3296
rect 23876 3232 23892 3296
rect 23956 3232 23972 3296
rect 24036 3232 24044 3296
rect 23644 2208 24044 3232
rect 23644 2144 23652 2208
rect 23716 2144 23732 2208
rect 23796 2144 23812 2208
rect 23876 2144 23892 2208
rect 23956 2144 23972 2208
rect 24036 2144 24044 2208
rect 23644 2128 24044 2144
<< via4 >>
rect 2986 24058 3222 24294
rect 2986 20160 3222 20294
rect 2986 20096 2992 20160
rect 2992 20096 3056 20160
rect 3056 20096 3072 20160
rect 3072 20096 3136 20160
rect 3136 20096 3152 20160
rect 3152 20096 3216 20160
rect 3216 20096 3222 20160
rect 2986 20058 3222 20096
rect 2986 16058 3222 16294
rect 2986 12058 3222 12294
rect 2986 8192 3222 8294
rect 2986 8128 2992 8192
rect 2992 8128 3056 8192
rect 3056 8128 3072 8192
rect 3072 8128 3136 8192
rect 3136 8128 3152 8192
rect 3152 8128 3216 8192
rect 3216 8128 3222 8192
rect 2986 8058 3222 8128
rect 2986 4058 3222 4294
rect 3726 24992 3732 25034
rect 3732 24992 3796 25034
rect 3796 24992 3812 25034
rect 3812 24992 3876 25034
rect 3876 24992 3892 25034
rect 3892 24992 3956 25034
rect 3956 24992 3962 25034
rect 3726 24798 3962 24992
rect 6986 24058 7222 24294
rect 3726 20798 3962 21034
rect 3726 16798 3962 17034
rect 3726 13024 3732 13034
rect 3732 13024 3796 13034
rect 3796 13024 3812 13034
rect 3812 13024 3876 13034
rect 3876 13024 3892 13034
rect 3892 13024 3956 13034
rect 3956 13024 3962 13034
rect 3726 12798 3962 13024
rect 3726 8798 3962 9034
rect 6986 20160 7222 20294
rect 6986 20096 6992 20160
rect 6992 20096 7056 20160
rect 7056 20096 7072 20160
rect 7072 20096 7136 20160
rect 7136 20096 7152 20160
rect 7152 20096 7216 20160
rect 7216 20096 7222 20160
rect 6986 20058 7222 20096
rect 6986 16058 7222 16294
rect 6986 12058 7222 12294
rect 6986 8192 7222 8294
rect 6986 8128 6992 8192
rect 6992 8128 7056 8192
rect 7056 8128 7072 8192
rect 7072 8128 7136 8192
rect 7136 8128 7152 8192
rect 7152 8128 7216 8192
rect 7216 8128 7222 8192
rect 6986 8058 7222 8128
rect 3726 4798 3962 5034
rect 6986 4058 7222 4294
rect 7726 24992 7732 25034
rect 7732 24992 7796 25034
rect 7796 24992 7812 25034
rect 7812 24992 7876 25034
rect 7876 24992 7892 25034
rect 7892 24992 7956 25034
rect 7956 24992 7962 25034
rect 7726 24798 7962 24992
rect 7726 20798 7962 21034
rect 7726 16798 7962 17034
rect 7726 13024 7732 13034
rect 7732 13024 7796 13034
rect 7796 13024 7812 13034
rect 7812 13024 7876 13034
rect 7876 13024 7892 13034
rect 7892 13024 7956 13034
rect 7956 13024 7962 13034
rect 7726 12798 7962 13024
rect 10986 24058 11222 24294
rect 10986 20160 11222 20294
rect 10986 20096 10992 20160
rect 10992 20096 11056 20160
rect 11056 20096 11072 20160
rect 11072 20096 11136 20160
rect 11136 20096 11152 20160
rect 11152 20096 11216 20160
rect 11216 20096 11222 20160
rect 10986 20058 11222 20096
rect 10986 16058 11222 16294
rect 10986 12058 11222 12294
rect 7726 8798 7962 9034
rect 7726 4798 7962 5034
rect 10986 8192 11222 8294
rect 10986 8128 10992 8192
rect 10992 8128 11056 8192
rect 11056 8128 11072 8192
rect 11072 8128 11136 8192
rect 11136 8128 11152 8192
rect 11152 8128 11216 8192
rect 11216 8128 11222 8192
rect 10986 8058 11222 8128
rect 10986 4058 11222 4294
rect 11726 24992 11732 25034
rect 11732 24992 11796 25034
rect 11796 24992 11812 25034
rect 11812 24992 11876 25034
rect 11876 24992 11892 25034
rect 11892 24992 11956 25034
rect 11956 24992 11962 25034
rect 11726 24798 11962 24992
rect 11726 20798 11962 21034
rect 14986 24058 15222 24294
rect 14986 20160 15222 20294
rect 14986 20096 14992 20160
rect 14992 20096 15056 20160
rect 15056 20096 15072 20160
rect 15072 20096 15136 20160
rect 15136 20096 15152 20160
rect 15152 20096 15216 20160
rect 15216 20096 15222 20160
rect 14986 20058 15222 20096
rect 11726 16798 11962 17034
rect 15726 24992 15732 25034
rect 15732 24992 15796 25034
rect 15796 24992 15812 25034
rect 15812 24992 15876 25034
rect 15876 24992 15892 25034
rect 15892 24992 15956 25034
rect 15956 24992 15962 25034
rect 15726 24798 15962 24992
rect 15726 20798 15962 21034
rect 15726 16798 15962 17034
rect 14986 16058 15222 16294
rect 11726 13024 11732 13034
rect 11732 13024 11796 13034
rect 11796 13024 11812 13034
rect 11812 13024 11876 13034
rect 11876 13024 11892 13034
rect 11892 13024 11956 13034
rect 11956 13024 11962 13034
rect 11726 12798 11962 13024
rect 11726 8798 11962 9034
rect 14986 12058 15222 12294
rect 11726 4798 11962 5034
rect 14986 8192 15222 8294
rect 14986 8128 14992 8192
rect 14992 8128 15056 8192
rect 15056 8128 15072 8192
rect 15072 8128 15136 8192
rect 15136 8128 15152 8192
rect 15152 8128 15216 8192
rect 15216 8128 15222 8192
rect 14986 8058 15222 8128
rect 14986 4058 15222 4294
rect 15726 13024 15732 13034
rect 15732 13024 15796 13034
rect 15796 13024 15812 13034
rect 15812 13024 15876 13034
rect 15876 13024 15892 13034
rect 15892 13024 15956 13034
rect 15956 13024 15962 13034
rect 15726 12798 15962 13024
rect 18986 24058 19222 24294
rect 19726 24992 19732 25034
rect 19732 24992 19796 25034
rect 19796 24992 19812 25034
rect 19812 24992 19876 25034
rect 19876 24992 19892 25034
rect 19892 24992 19956 25034
rect 19956 24992 19962 25034
rect 19726 24798 19962 24992
rect 18986 20160 19222 20294
rect 18986 20096 18992 20160
rect 18992 20096 19056 20160
rect 19056 20096 19072 20160
rect 19072 20096 19136 20160
rect 19136 20096 19152 20160
rect 19152 20096 19216 20160
rect 19216 20096 19222 20160
rect 18986 20058 19222 20096
rect 15726 8798 15962 9034
rect 18986 16058 19222 16294
rect 19726 20798 19962 21034
rect 19726 16798 19962 17034
rect 18986 12058 19222 12294
rect 18986 8192 19222 8294
rect 18986 8128 18992 8192
rect 18992 8128 19056 8192
rect 19056 8128 19072 8192
rect 19072 8128 19136 8192
rect 19136 8128 19152 8192
rect 19152 8128 19216 8192
rect 19216 8128 19222 8192
rect 18986 8058 19222 8128
rect 15726 4798 15962 5034
rect 18986 4058 19222 4294
rect 19726 13024 19732 13034
rect 19732 13024 19796 13034
rect 19796 13024 19812 13034
rect 19812 13024 19876 13034
rect 19876 13024 19892 13034
rect 19892 13024 19956 13034
rect 19956 13024 19962 13034
rect 19726 12798 19962 13024
rect 19726 8798 19962 9034
rect 19726 4798 19962 5034
rect 22986 24058 23222 24294
rect 22986 20160 23222 20294
rect 22986 20096 22992 20160
rect 22992 20096 23056 20160
rect 23056 20096 23072 20160
rect 23072 20096 23136 20160
rect 23136 20096 23152 20160
rect 23152 20096 23216 20160
rect 23216 20096 23222 20160
rect 22986 20058 23222 20096
rect 22986 16058 23222 16294
rect 22986 12058 23222 12294
rect 22986 8192 23222 8294
rect 22986 8128 22992 8192
rect 22992 8128 23056 8192
rect 23056 8128 23072 8192
rect 23072 8128 23136 8192
rect 23136 8128 23152 8192
rect 23152 8128 23216 8192
rect 23216 8128 23222 8192
rect 22986 8058 23222 8128
rect 22986 4058 23222 4294
rect 23726 24992 23732 25034
rect 23732 24992 23796 25034
rect 23796 24992 23812 25034
rect 23812 24992 23876 25034
rect 23876 24992 23892 25034
rect 23892 24992 23956 25034
rect 23956 24992 23962 25034
rect 23726 24798 23962 24992
rect 23726 20798 23962 21034
rect 23726 16798 23962 17034
rect 23726 13024 23732 13034
rect 23732 13024 23796 13034
rect 23796 13024 23812 13034
rect 23812 13024 23876 13034
rect 23876 13024 23892 13034
rect 23892 13024 23956 13034
rect 23956 13024 23962 13034
rect 23726 12798 23962 13024
rect 23726 8798 23962 9034
rect 23726 4798 23962 5034
<< metal5 >>
rect 1056 25034 26912 25116
rect 1056 24798 3726 25034
rect 3962 24798 7726 25034
rect 7962 24798 11726 25034
rect 11962 24798 15726 25034
rect 15962 24798 19726 25034
rect 19962 24798 23726 25034
rect 23962 24798 26912 25034
rect 1056 24716 26912 24798
rect 1056 24294 26912 24376
rect 1056 24058 2986 24294
rect 3222 24058 6986 24294
rect 7222 24058 10986 24294
rect 11222 24058 14986 24294
rect 15222 24058 18986 24294
rect 19222 24058 22986 24294
rect 23222 24058 26912 24294
rect 1056 23976 26912 24058
rect 1056 21034 26912 21116
rect 1056 20798 3726 21034
rect 3962 20798 7726 21034
rect 7962 20798 11726 21034
rect 11962 20798 15726 21034
rect 15962 20798 19726 21034
rect 19962 20798 23726 21034
rect 23962 20798 26912 21034
rect 1056 20716 26912 20798
rect 1056 20294 26912 20376
rect 1056 20058 2986 20294
rect 3222 20058 6986 20294
rect 7222 20058 10986 20294
rect 11222 20058 14986 20294
rect 15222 20058 18986 20294
rect 19222 20058 22986 20294
rect 23222 20058 26912 20294
rect 1056 19976 26912 20058
rect 1056 17034 26912 17116
rect 1056 16798 3726 17034
rect 3962 16798 7726 17034
rect 7962 16798 11726 17034
rect 11962 16798 15726 17034
rect 15962 16798 19726 17034
rect 19962 16798 23726 17034
rect 23962 16798 26912 17034
rect 1056 16716 26912 16798
rect 1056 16294 26912 16376
rect 1056 16058 2986 16294
rect 3222 16058 6986 16294
rect 7222 16058 10986 16294
rect 11222 16058 14986 16294
rect 15222 16058 18986 16294
rect 19222 16058 22986 16294
rect 23222 16058 26912 16294
rect 1056 15976 26912 16058
rect 1056 13034 26912 13116
rect 1056 12798 3726 13034
rect 3962 12798 7726 13034
rect 7962 12798 11726 13034
rect 11962 12798 15726 13034
rect 15962 12798 19726 13034
rect 19962 12798 23726 13034
rect 23962 12798 26912 13034
rect 1056 12716 26912 12798
rect 1056 12294 26912 12376
rect 1056 12058 2986 12294
rect 3222 12058 6986 12294
rect 7222 12058 10986 12294
rect 11222 12058 14986 12294
rect 15222 12058 18986 12294
rect 19222 12058 22986 12294
rect 23222 12058 26912 12294
rect 1056 11976 26912 12058
rect 1056 9034 26912 9116
rect 1056 8798 3726 9034
rect 3962 8798 7726 9034
rect 7962 8798 11726 9034
rect 11962 8798 15726 9034
rect 15962 8798 19726 9034
rect 19962 8798 23726 9034
rect 23962 8798 26912 9034
rect 1056 8716 26912 8798
rect 1056 8294 26912 8376
rect 1056 8058 2986 8294
rect 3222 8058 6986 8294
rect 7222 8058 10986 8294
rect 11222 8058 14986 8294
rect 15222 8058 18986 8294
rect 19222 8058 22986 8294
rect 23222 8058 26912 8294
rect 1056 7976 26912 8058
rect 1056 5034 26912 5116
rect 1056 4798 3726 5034
rect 3962 4798 7726 5034
rect 7962 4798 11726 5034
rect 11962 4798 15726 5034
rect 15962 4798 19726 5034
rect 19962 4798 23726 5034
rect 23962 4798 26912 5034
rect 1056 4716 26912 4798
rect 1056 4294 26912 4376
rect 1056 4058 2986 4294
rect 3222 4058 6986 4294
rect 7222 4058 10986 4294
rect 11222 4058 14986 4294
rect 15222 4058 18986 4294
rect 19222 4058 22986 4294
rect 23222 4058 26912 4294
rect 1056 3976 26912 4058
use sky130_fd_sc_hd__buf_2  _0547_
timestamp 0
transform -1 0 24288 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0548_
timestamp 0
transform -1 0 23920 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0549_
timestamp 0
transform 1 0 23184 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0550_
timestamp 0
transform 1 0 25668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0551_
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0552_
timestamp 0
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0553_
timestamp 0
transform -1 0 22448 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0554_
timestamp 0
transform 1 0 24564 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0555_
timestamp 0
transform 1 0 25576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0556_
timestamp 0
transform 1 0 25208 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0557_
timestamp 0
transform -1 0 25576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 0
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0559_
timestamp 0
transform -1 0 25852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0560_
timestamp 0
transform -1 0 25116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 0
transform -1 0 24748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0562_
timestamp 0
transform 1 0 23920 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0563_
timestamp 0
transform 1 0 23092 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0564_
timestamp 0
transform 1 0 22908 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0565_
timestamp 0
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0566_
timestamp 0
transform -1 0 23368 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0567_
timestamp 0
transform -1 0 25484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0568_
timestamp 0
transform -1 0 25668 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0569_
timestamp 0
transform 1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0570_
timestamp 0
transform -1 0 18216 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0571_
timestamp 0
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0572_
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0573_
timestamp 0
transform 1 0 20792 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0574_
timestamp 0
transform -1 0 23276 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0575_
timestamp 0
transform 1 0 21988 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 0
transform -1 0 24472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0578_
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 0
transform 1 0 23736 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0580_
timestamp 0
transform -1 0 25576 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0581_
timestamp 0
transform 1 0 24840 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 0
transform -1 0 24748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 0
transform -1 0 21712 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 0
transform 1 0 20792 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 0
transform 1 0 20608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0586_
timestamp 0
transform 1 0 22172 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0587_
timestamp 0
transform 1 0 21712 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0588_
timestamp 0
transform 1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 0
transform 1 0 25208 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0591_
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0592_
timestamp 0
transform 1 0 23552 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0593_
timestamp 0
transform -1 0 25300 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 0
transform -1 0 25208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 0
transform -1 0 25576 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0596_
timestamp 0
transform -1 0 25300 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0597_
timestamp 0
transform 1 0 22356 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0598_
timestamp 0
transform -1 0 26128 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0599_
timestamp 0
transform 1 0 24288 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0600_
timestamp 0
transform 1 0 23552 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _0601_
timestamp 0
transform 1 0 24932 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 0
transform -1 0 24748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 0
transform 1 0 23920 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0604_
timestamp 0
transform 1 0 23552 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0605_
timestamp 0
transform 1 0 24104 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0606_
timestamp 0
transform 1 0 21528 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0607_
timestamp 0
transform -1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0608_
timestamp 0
transform 1 0 19044 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0609_
timestamp 0
transform 1 0 19872 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0610_
timestamp 0
transform 1 0 20424 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0611_
timestamp 0
transform 1 0 20240 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0612_
timestamp 0
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0613_
timestamp 0
transform -1 0 21344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0614_
timestamp 0
transform 1 0 21528 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0615_
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0616_
timestamp 0
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0617_
timestamp 0
transform -1 0 20148 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0618_
timestamp 0
transform 1 0 22264 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 0
transform 1 0 23276 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 0
transform -1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0621_
timestamp 0
transform 1 0 21988 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0622_
timestamp 0
transform 1 0 20884 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 0
transform -1 0 22816 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 0
transform -1 0 22448 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0625_
timestamp 0
transform 1 0 20240 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0626_
timestamp 0
transform 1 0 20424 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 0
transform -1 0 24012 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0628_
timestamp 0
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 0
transform 1 0 22080 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 0
transform -1 0 21528 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 0
transform -1 0 22080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0632_
timestamp 0
transform -1 0 20608 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0633_
timestamp 0
transform 1 0 19688 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0634_
timestamp 0
transform 1 0 19596 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0635_
timestamp 0
transform 1 0 20148 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0636_
timestamp 0
transform -1 0 20148 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0637_
timestamp 0
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0638_
timestamp 0
transform -1 0 19504 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0639_
timestamp 0
transform -1 0 21436 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0640_
timestamp 0
transform 1 0 15916 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0641_
timestamp 0
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_4  _0642_
timestamp 0
transform 1 0 17480 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__and3b_4  _0643_
timestamp 0
transform -1 0 20240 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0644_
timestamp 0
transform -1 0 19320 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_4  _0645_
timestamp 0
transform -1 0 17940 0 1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__a22o_1  _0646_
timestamp 0
transform 1 0 12972 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_4  _0647_
timestamp 0
transform -1 0 20424 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0648_
timestamp 0
transform -1 0 14720 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0649_
timestamp 0
transform -1 0 18124 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0650_
timestamp 0
transform 1 0 13892 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0651_
timestamp 0
transform 1 0 16652 0 1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__nor4b_4  _0652_
timestamp 0
transform -1 0 20056 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__a22o_1  _0653_
timestamp 0
transform 1 0 13156 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0654_
timestamp 0
transform 1 0 18124 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and4bb_4  _0655_
timestamp 0
transform 1 0 17940 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and4b_4  _0656_
timestamp 0
transform -1 0 19044 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__and4bb_4  _0657_
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0658_
timestamp 0
transform -1 0 14536 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0659_
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_4  _0660_
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__nor4b_4  _0661_
timestamp 0
transform -1 0 17940 0 1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__and4bb_4  _0662_
timestamp 0
transform 1 0 17940 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and4bb_4  _0663_
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0664_
timestamp 0
transform 1 0 12696 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0665_
timestamp 0
transform 1 0 13800 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0666_
timestamp 0
transform 1 0 14168 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0667_
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0668_
timestamp 0
transform -1 0 20608 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0669_
timestamp 0
transform -1 0 14536 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0670_
timestamp 0
transform -1 0 13984 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0671_
timestamp 0
transform 1 0 16744 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0672_
timestamp 0
transform -1 0 17756 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0673_
timestamp 0
transform 1 0 16284 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0674_
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0675_
timestamp 0
transform 1 0 15916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0676_
timestamp 0
transform -1 0 18124 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0677_
timestamp 0
transform -1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0678_
timestamp 0
transform 1 0 16928 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0679_
timestamp 0
transform -1 0 17572 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0680_
timestamp 0
transform 1 0 16836 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0681_
timestamp 0
transform 1 0 17480 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0682_
timestamp 0
transform 1 0 13248 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0683_
timestamp 0
transform 1 0 12972 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0684_
timestamp 0
transform -1 0 11040 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0685_
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0686_
timestamp 0
transform 1 0 7820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0687_
timestamp 0
transform 1 0 6348 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0688_
timestamp 0
transform 1 0 6716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0689_
timestamp 0
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0690_
timestamp 0
transform -1 0 12236 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0691_
timestamp 0
transform 1 0 12144 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0692_
timestamp 0
transform -1 0 12144 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0693_
timestamp 0
transform 1 0 10856 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0694_
timestamp 0
transform 1 0 10488 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 0
transform 1 0 4140 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0696_
timestamp 0
transform -1 0 7360 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0697_
timestamp 0
transform 1 0 3772 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0698_
timestamp 0
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0699_
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0700_
timestamp 0
transform 1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0701_
timestamp 0
transform 1 0 5796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0702_
timestamp 0
transform 1 0 10120 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0703_
timestamp 0
transform -1 0 9568 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0704_
timestamp 0
transform 1 0 9752 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0705_
timestamp 0
transform 1 0 4784 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0706_
timestamp 0
transform -1 0 9660 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 0
transform -1 0 9844 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0708_
timestamp 0
transform 1 0 8096 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0709_
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0710_
timestamp 0
transform 1 0 7636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0711_
timestamp 0
transform -1 0 11316 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0712_
timestamp 0
transform 1 0 8096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0713_
timestamp 0
transform 1 0 8924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0714_
timestamp 0
transform -1 0 10120 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0715_
timestamp 0
transform -1 0 9568 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0716_
timestamp 0
transform 1 0 10672 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0717_
timestamp 0
transform 1 0 9936 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0718_
timestamp 0
transform 1 0 10396 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 0
transform 1 0 5152 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0720_
timestamp 0
transform 1 0 6256 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0721_
timestamp 0
transform -1 0 5244 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0722_
timestamp 0
transform 1 0 4232 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0723_
timestamp 0
transform 1 0 3772 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0724_
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0725_
timestamp 0
transform -1 0 6256 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0726_
timestamp 0
transform -1 0 10120 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0727_
timestamp 0
transform -1 0 10028 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0728_
timestamp 0
transform 1 0 10028 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0729_
timestamp 0
transform 1 0 10396 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0730_
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0731_
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0732_
timestamp 0
transform -1 0 8464 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0733_
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0734_
timestamp 0
transform 1 0 4600 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0735_
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0736_
timestamp 0
transform 1 0 4784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0737_
timestamp 0
transform 1 0 5612 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0738_
timestamp 0
transform 1 0 10396 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0739_
timestamp 0
transform -1 0 10120 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0740_
timestamp 0
transform 1 0 10304 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp 0
transform 1 0 15364 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0742_
timestamp 0
transform -1 0 16836 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0743_
timestamp 0
transform 1 0 19596 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0744_
timestamp 0
transform 1 0 18400 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0745_
timestamp 0
transform 1 0 18492 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0746_
timestamp 0
transform -1 0 19044 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0747_
timestamp 0
transform 1 0 15732 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0748_
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0749_
timestamp 0
transform 1 0 20056 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0750_
timestamp 0
transform -1 0 19596 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0751_
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0752_
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0753_
timestamp 0
transform -1 0 21712 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0755_
timestamp 0
transform 1 0 22816 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0756_
timestamp 0
transform -1 0 22724 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 0
transform -1 0 21712 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 0
transform -1 0 26128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 0
transform 1 0 26220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 0
transform -1 0 23736 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 0
transform -1 0 23092 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 0
transform 1 0 22080 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 0
transform 1 0 26128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 0
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 0
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 0
transform -1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0767_
timestamp 0
transform -1 0 21160 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 0
transform 1 0 20240 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 0
transform -1 0 12328 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 0
transform -1 0 12236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 0
transform -1 0 11776 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 0
transform -1 0 11408 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 0
transform -1 0 12512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 0
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 0
transform -1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 0
transform 1 0 17388 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 0
transform -1 0 20884 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 0
transform -1 0 22264 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 0
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 0
transform -1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0781_
timestamp 0
transform -1 0 21712 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0782_
timestamp 0
transform 1 0 23552 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 0
transform -1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 0
transform -1 0 23092 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 0
transform 1 0 26220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 0
transform -1 0 23276 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 0
transform -1 0 23552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 0
transform 1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 0
transform 1 0 25024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 0
transform 1 0 24104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 0
transform -1 0 23184 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 0
transform -1 0 22080 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 0
transform 1 0 24656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 0
transform 1 0 23184 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 0
transform -1 0 25944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 0
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 0
transform 1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 0
transform 1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 0
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 0
transform 1 0 25484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 0
transform -1 0 25484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 0
transform -1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 0
transform 1 0 22448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0806_
timestamp 0
transform -1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _0807_
timestamp 0
transform -1 0 23276 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0808_
timestamp 0
transform -1 0 18584 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_4  _0809_
timestamp 0
transform -1 0 21344 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0811_
timestamp 0
transform -1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0812_
timestamp 0
transform -1 0 4140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 0
transform -1 0 9292 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0814_
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0815_
timestamp 0
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0817_
timestamp 0
transform 1 0 7084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0818_
timestamp 0
transform -1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp 0
transform 1 0 7912 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 0
transform 1 0 7636 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0821_
timestamp 0
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 0
transform 1 0 9108 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0823_
timestamp 0
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0824_
timestamp 0
transform -1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 0
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0827_
timestamp 0
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 0
transform 1 0 17388 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0829_
timestamp 0
transform -1 0 17480 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0830_
timestamp 0
transform -1 0 13708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 0
transform 1 0 12972 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 0
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0833_
timestamp 0
transform -1 0 20700 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_4  _0834_
timestamp 0
transform -1 0 20700 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 0
transform 1 0 14536 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 0
transform 1 0 14260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp 0
transform 1 0 2760 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0838_
timestamp 0
transform 1 0 2300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0839_
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0840_
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0841_
timestamp 0
transform 1 0 7176 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0842_
timestamp 0
transform -1 0 6624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0843_
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 0
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 0
transform 1 0 9476 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 0
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0847_
timestamp 0
transform -1 0 16836 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0848_
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 0
transform 1 0 13340 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0850_
timestamp 0
transform -1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0851_
timestamp 0
transform -1 0 22908 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_4  _0852_
timestamp 0
transform -1 0 21160 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 0
transform -1 0 19780 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0854_
timestamp 0
transform -1 0 20056 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 0
transform -1 0 6256 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0856_
timestamp 0
transform -1 0 6440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 0
transform -1 0 8188 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0858_
timestamp 0
transform 1 0 8188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 0
transform 1 0 4048 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 0
transform 1 0 3036 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0862_
timestamp 0
transform -1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp 0
transform 1 0 6256 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0864_
timestamp 0
transform -1 0 6164 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0865_
timestamp 0
transform -1 0 18860 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0866_
timestamp 0
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 0
transform 1 0 12328 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0868_
timestamp 0
transform 1 0 12052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0869_
timestamp 0
transform -1 0 21620 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_4  _0870_
timestamp 0
transform -1 0 22172 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0871_
timestamp 0
transform -1 0 19228 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 0
transform -1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 0
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0874_
timestamp 0
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0875_
timestamp 0
transform 1 0 4876 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0876_
timestamp 0
transform 1 0 4692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0877_
timestamp 0
transform 1 0 4876 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp 0
transform 1 0 7268 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0880_
timestamp 0
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0881_
timestamp 0
transform 1 0 6992 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0882_
timestamp 0
transform 1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0883_
timestamp 0
transform 1 0 15640 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 0
transform 1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0885_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 0
transform -1 0 13616 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _0887_
timestamp 0
transform 1 0 19964 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_4  _0888_
timestamp 0
transform -1 0 20148 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0889_
timestamp 0
transform 1 0 14444 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0890_
timestamp 0
transform -1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0891_
timestamp 0
transform 1 0 3496 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0892_
timestamp 0
transform -1 0 2024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 0
transform 1 0 5428 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0894_
timestamp 0
transform 1 0 5244 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0895_
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0896_
timestamp 0
transform 1 0 4600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0897_
timestamp 0
transform 1 0 10672 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 0
transform -1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0900_
timestamp 0
transform -1 0 6624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0901_
timestamp 0
transform 1 0 14628 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0902_
timestamp 0
transform 1 0 14352 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0903_
timestamp 0
transform 1 0 12236 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 0
transform -1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _0905_
timestamp 0
transform -1 0 20700 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 0
transform 1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 0
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0908_
timestamp 0
transform 1 0 2668 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 0
transform 1 0 2300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 0
transform 1 0 4048 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 0
transform 1 0 3864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0912_
timestamp 0
transform 1 0 5060 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 0
transform 1 0 4784 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 0
transform 1 0 3036 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 0
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp 0
transform 1 0 9568 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 0
transform -1 0 9292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 0
transform 1 0 14904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 0
transform 1 0 14352 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 0
transform -1 0 12880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0922_
timestamp 0
transform -1 0 23828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0923_
timestamp 0
transform -1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_4  _0924_
timestamp 0
transform -1 0 19872 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0925_
timestamp 0
transform 1 0 14352 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0926_
timestamp 0
transform -1 0 13616 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0927_
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0928_
timestamp 0
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 0
transform 1 0 3128 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0930_
timestamp 0
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0931_
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0932_
timestamp 0
transform 1 0 7820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0933_
timestamp 0
transform 1 0 2024 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0934_
timestamp 0
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp 0
transform 1 0 6992 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 0
transform -1 0 6256 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0937_
timestamp 0
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0938_
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 0
transform 1 0 13064 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0940_
timestamp 0
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _0941_
timestamp 0
transform -1 0 20700 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 0
transform 1 0 18952 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 0
transform -1 0 19044 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp 0
transform 1 0 3956 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 0
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 0
transform 1 0 3772 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 0
transform 1 0 7820 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 0
transform 1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 0
transform 1 0 4048 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 0
transform 1 0 11776 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0953_
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 0
transform -1 0 18860 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 0
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 0
transform 1 0 14168 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 0
transform 1 0 13340 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _0958_
timestamp 0
transform -1 0 19136 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_4  _0959_
timestamp 0
transform -1 0 19688 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 0
transform -1 0 14444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0962_
timestamp 0
transform 1 0 2760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 0
transform 1 0 2392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp 0
transform 1 0 2852 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 0
transform 1 0 2392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp 0
transform 1 0 7912 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 0
transform 1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 0
transform 1 0 2208 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0969_
timestamp 0
transform -1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 0
transform 1 0 11960 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 0
transform -1 0 11500 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0972_
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 0
transform -1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0974_
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0975_
timestamp 0
transform 1 0 13064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _0976_
timestamp 0
transform -1 0 19688 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0977_
timestamp 0
transform 1 0 15732 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 0
transform 1 0 15088 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp 0
transform -1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 0
transform -1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 0
transform 1 0 5888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0983_
timestamp 0
transform -1 0 8372 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 0
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0985_
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 0
transform 1 0 6348 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0987_
timestamp 0
transform 1 0 7912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 0
transform 1 0 6716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0989_
timestamp 0
transform 1 0 15548 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 0
transform 1 0 15272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp 0
transform 1 0 13340 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 0
transform 1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _0993_
timestamp 0
transform -1 0 19136 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 0
transform 1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 0
transform 1 0 4324 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 0
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 0
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 0
transform 1 0 2852 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 0
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 0
transform 1 0 5428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 0
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 0
transform 1 0 15548 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 0
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 0
transform -1 0 12144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _1010_
timestamp 0
transform -1 0 20700 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 0
transform 1 0 17940 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 0
transform -1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1013_
timestamp 0
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1015_
timestamp 0
transform -1 0 5428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 0
transform 1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 0
transform 1 0 7452 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 0
transform -1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 0
transform 1 0 4324 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 0
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 0
transform 1 0 12144 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 0
transform -1 0 11776 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1023_
timestamp 0
transform 1 0 15916 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 0
transform 1 0 15548 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 0
transform 1 0 12972 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 0
transform 1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1027_
timestamp 0
transform 1 0 20700 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_4  _1028_
timestamp 0
transform 1 0 20700 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 0
transform 1 0 17480 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 0
transform 1 0 16744 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1031_
timestamp 0
transform 1 0 3772 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 0
transform 1 0 2760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1033_
timestamp 0
transform 1 0 2944 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 0
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1035_
timestamp 0
transform -1 0 9476 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 0
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1037_
timestamp 0
transform 1 0 4968 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 0
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1039_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 0
transform 1 0 5888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1041_
timestamp 0
transform 1 0 15640 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 0
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1043_
timestamp 0
transform 1 0 13064 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1044_
timestamp 0
transform 1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _1045_
timestamp 0
transform -1 0 21160 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1046_
timestamp 0
transform 1 0 16744 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 0
transform 1 0 10488 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 0
transform 1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 0
transform 1 0 9292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 0
transform 1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1052_
timestamp 0
transform -1 0 10672 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 0
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1054_
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 0
transform -1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1056_
timestamp 0
transform 1 0 10212 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 0
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1058_
timestamp 0
transform -1 0 18768 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1059_
timestamp 0
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1060_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 0
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _1062_
timestamp 0
transform -1 0 19964 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1063_
timestamp 0
transform 1 0 18124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 0
transform -1 0 16744 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1065_
timestamp 0
transform 1 0 6532 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1067_
timestamp 0
transform 1 0 9016 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 0
transform -1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1069_
timestamp 0
transform 1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 0
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1071_
timestamp 0
transform 1 0 6624 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 0
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1073_
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 0
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1075_
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 0
transform -1 0 16376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1077_
timestamp 0
transform 1 0 13340 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 0
transform 1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_4  _1079_
timestamp 0
transform -1 0 22172 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1080_
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 0
transform -1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1082_
timestamp 0
transform -1 0 10948 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1083_
timestamp 0
transform -1 0 11224 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1084_
timestamp 0
transform 1 0 9384 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1085_
timestamp 0
transform 1 0 9292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1086_
timestamp 0
transform 1 0 9844 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1087_
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1088_
timestamp 0
transform 1 0 10488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 0
transform -1 0 9292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1090_
timestamp 0
transform 1 0 13156 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1091_
timestamp 0
transform -1 0 11408 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1092_
timestamp 0
transform -1 0 17940 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1093_
timestamp 0
transform -1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1094_
timestamp 0
transform 1 0 13248 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1095_
timestamp 0
transform -1 0 12052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 0
transform 1 0 20700 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 0
transform -1 0 26404 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1099_
timestamp 0
transform 1 0 21620 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 0
transform -1 0 23644 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 0
transform -1 0 23644 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 0
transform 1 0 24656 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 0
transform -1 0 26588 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 0
transform 1 0 22172 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 0
transform 1 0 10212 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 0
transform 1 0 10120 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 0
transform -1 0 11408 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 0
transform 1 0 9568 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 0
transform 1 0 10396 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 0
transform 1 0 15732 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 0
transform 1 0 12972 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1114_
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1115_
timestamp 0
transform -1 0 19780 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 0
transform 1 0 20148 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 0
transform -1 0 21712 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 0
transform 1 0 19872 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 0
transform 1 0 24380 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 0
transform 1 0 21160 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 0
transform 1 0 21436 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 0
transform 1 0 24748 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 0
transform -1 0 26404 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 0
transform 1 0 21988 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 0
transform -1 0 22356 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 0
transform 1 0 23644 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 0
transform 1 0 22448 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 0
transform 1 0 23460 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1132_
timestamp 0
transform 1 0 22172 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1133_
timestamp 0
transform 1 0 24472 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 0
transform 1 0 23092 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1135_
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1136_
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 0
transform 1 0 19872 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 0
transform 1 0 23368 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1140_
timestamp 0
transform 1 0 20884 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1141_
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 0
transform 1 0 18768 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 0
transform 1 0 7360 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 0
transform 1 0 6992 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 0
transform 1 0 7360 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 0
transform 1 0 11040 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 0
transform -1 0 19044 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 0
transform 1 0 12420 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 0
transform 1 0 13616 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 0
transform 1 0 1932 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 0
transform 1 0 2024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 0
transform 1 0 6624 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 0
transform 1 0 1932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 0
transform 1 0 15088 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 0
transform 1 0 11868 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 0
transform -1 0 20792 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 0
transform -1 0 8464 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 0
transform 1 0 2576 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 0
transform 1 0 1932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 0
transform -1 0 19320 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 0
transform 1 0 11684 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 0
transform -1 0 20700 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 0
transform 1 0 4140 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 0
transform 1 0 4232 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 0
transform 1 0 4048 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 0
transform 1 0 6716 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 0
transform 1 0 6440 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 0
transform 1 0 14168 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 0
transform 1 0 13616 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 0
transform 1 0 14444 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 0
transform 1 0 2024 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 0
transform 1 0 4324 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1178_
timestamp 0
transform 1 0 9016 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 0
transform 1 0 6716 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 0
transform 1 0 11776 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 0
transform 1 0 17664 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 0
transform 1 0 1840 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 0
transform 1 0 4416 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 0
transform 1 0 1564 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 0
transform 1 0 9660 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 0
transform 1 0 14260 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 0
transform 1 0 12880 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 0
transform 1 0 1472 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 0
transform 1 0 1656 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 0
transform 1 0 7544 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 0
transform 1 0 1472 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 0
transform 1 0 6440 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 0
transform 1 0 14904 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 0
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1200_
timestamp 0
transform 1 0 2208 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 0
transform 1 0 3496 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 0
transform 1 0 11040 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1204_
timestamp 0
transform -1 0 19136 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 0
transform 1 0 12512 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 0
transform 1 0 14260 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 0
transform 1 0 1932 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1208_
timestamp 0
transform 1 0 1932 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1209_
timestamp 0
transform 1 0 6440 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1210_
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1211_
timestamp 0
transform 1 0 11684 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1212_
timestamp 0
transform 1 0 15088 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp 0
transform 1 0 12696 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp 0
transform 1 0 14720 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp 0
transform -1 0 12880 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1216_
timestamp 0
transform 1 0 5336 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp 0
transform -1 0 8556 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1218_
timestamp 0
transform 1 0 5888 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1219_
timestamp 0
transform 1 0 6624 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1220_
timestamp 0
transform 1 0 14904 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1221_
timestamp 0
transform 1 0 12512 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1222_
timestamp 0
transform 1 0 15088 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1223_
timestamp 0
transform 1 0 1840 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1224_
timestamp 0
transform 1 0 2852 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1225_
timestamp 0
transform 1 0 6808 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1226_
timestamp 0
transform 1 0 1932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1227_
timestamp 0
transform 1 0 3956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1228_
timestamp 0
transform 1 0 14812 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1229_
timestamp 0
transform 1 0 11868 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1230_
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1231_
timestamp 0
transform 1 0 8464 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1232_
timestamp 0
transform 1 0 3956 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 0
transform 1 0 6900 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 0
transform 1 0 11776 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 0
transform 1 0 14996 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 0
transform 1 0 2300 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 0
transform 1 0 1472 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 0
transform 1 0 9200 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 0
transform 1 0 5520 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 0
transform 1 0 14996 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 0
transform 1 0 12512 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 0
transform 1 0 15272 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 0
transform 1 0 9016 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 0
transform -1 0 10948 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 0
transform 1 0 9384 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 0
transform 1 0 9660 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 0
transform -1 0 18492 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 0
transform 1 0 13064 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 0
transform 1 0 17020 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 0
transform 1 0 8464 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 0
transform 1 0 9200 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 0
transform 1 0 5152 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 0
transform 1 0 16468 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 0
transform 1 0 12144 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 0
transform -1 0 20700 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 0
transform -1 0 11408 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 0
transform 1 0 8924 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 0
transform 1 0 9476 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 0
transform 1 0 9292 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 0
transform 1 0 11868 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 0
transform -1 0 18400 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 0
transform 1 0 12052 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform -1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_rd_clk
timestamp 0
transform -1 0 19872 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wr_clk
timestamp 0
transform 1 0 13984 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_rd_clk
timestamp 0
transform -1 0 18492 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_rd_clk
timestamp 0
transform 1 0 20240 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_wr_clk
timestamp 0
transform 1 0 5152 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_wr_clk
timestamp 0
transform 1 0 4968 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_wr_clk
timestamp 0
transform -1 0 10672 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_wr_clk
timestamp 0
transform 1 0 9476 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_wr_clk
timestamp 0
transform -1 0 5520 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_wr_clk
timestamp 0
transform -1 0 6072 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_wr_clk
timestamp 0
transform 1 0 10396 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_wr_clk
timestamp 0
transform 1 0 10396 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_wr_clk
timestamp 0
transform -1 0 15916 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_wr_clk
timestamp 0
transform 1 0 14536 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_wr_clk
timestamp 0
transform 1 0 22172 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_wr_clk
timestamp 0
transform 1 0 20700 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_wr_clk
timestamp 0
transform -1 0 17664 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_wr_clk
timestamp 0
transform -1 0 17480 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_wr_clk
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_wr_clk
timestamp 0
transform 1 0 22540 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  clkload0
timestamp 0
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload2
timestamp 0
transform 1 0 9016 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload3
timestamp 0
transform 1 0 8832 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload4
timestamp 0
transform 1 0 4508 0 1 19584
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  clkload5
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload6
timestamp 0
transform 1 0 10396 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload7
timestamp 0
transform 1 0 14444 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload8
timestamp 0
transform 1 0 14444 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload9
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload10
timestamp 0
transform -1 0 21344 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload11
timestamp 0
transform 1 0 15916 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload12
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload13
timestamp 0
transform 1 0 21436 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload14
timestamp 0
transform 1 0 21068 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload15
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_65
timestamp 0
transform 1 0 7084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_73
timestamp 0
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_95
timestamp 0
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_107
timestamp 0
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 0
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_161
timestamp 0
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_177
timestamp 0
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_189
timestamp 0
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 0
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 0
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_78
timestamp 0
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_86
timestamp 0
transform 1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_104
timestamp 0
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_142
timestamp 0
transform 1 0 14168 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_154
timestamp 0
transform 1 0 15272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_158
timestamp 0
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_162
timestamp 0
transform 1 0 16008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 0
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_189
timestamp 0
transform 1 0 18492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_201
timestamp 0
transform 1 0 19596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_213
timestamp 0
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_221
timestamp 0
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_231
timestamp 0
transform 1 0 22356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_235
timestamp 0
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_259
timestamp 0
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_271
timestamp 0
transform 1 0 26036 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_40
timestamp 0
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_60
timestamp 0
transform 1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_78
timestamp 0
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_104
timestamp 0
transform 1 0 10672 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_116
timestamp 0
transform 1 0 11776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_136
timestamp 0
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_150
timestamp 0
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_213
timestamp 0
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_244
timestamp 0
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_256
timestamp 0
transform 1 0 24656 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_261
timestamp 0
transform 1 0 25116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_273
timestamp 0
transform 1 0 26220 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_48
timestamp 0
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 0
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_79
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 0
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_121
timestamp 0
transform 1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_126
timestamp 0
transform 1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_146
timestamp 0
transform 1 0 14536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_185
timestamp 0
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_212
timestamp 0
transform 1 0 20608 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_248
timestamp 0
transform 1 0 23920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_272
timestamp 0
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_276
timestamp 0
transform 1 0 26496 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_32
timestamp 0
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_36
timestamp 0
transform 1 0 4416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_40
timestamp 0
transform 1 0 4784 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_46
timestamp 0
transform 1 0 5336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_54
timestamp 0
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_64
timestamp 0
transform 1 0 6992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_68
timestamp 0
transform 1 0 7360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_78
timestamp 0
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_111
timestamp 0
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_123
timestamp 0
transform 1 0 12420 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_149
timestamp 0
transform 1 0 14812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_161
timestamp 0
transform 1 0 15916 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_218
timestamp 0
transform 1 0 21160 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_235
timestamp 0
transform 1 0 22724 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_243
timestamp 0
transform 1 0 23460 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_247
timestamp 0
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_256
timestamp 0
transform 1 0 24656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_268
timestamp 0
transform 1 0 25760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_276
timestamp 0
transform 1 0 26496 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_31
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 0
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_79
timestamp 0
transform 1 0 8372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_91
timestamp 0
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_101
timestamp 0
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 0
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_132
timestamp 0
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_172
timestamp 0
transform 1 0 16928 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_218
timestamp 0
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 0
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 0
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 0
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_273
timestamp 0
transform 1 0 26220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 0
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_64
timestamp 0
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_80
timestamp 0
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_93
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_104
timestamp 0
transform 1 0 10672 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_116
timestamp 0
transform 1 0 11776 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_120
timestamp 0
transform 1 0 12144 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_132
timestamp 0
transform 1 0 13248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 0
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_150
timestamp 0
transform 1 0 14904 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_171
timestamp 0
transform 1 0 16836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_179
timestamp 0
transform 1 0 17572 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_237
timestamp 0
transform 1 0 22908 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_245
timestamp 0
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_271
timestamp 0
transform 1 0 26036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_34
timestamp 0
transform 1 0 4232 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_44
timestamp 0
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_82
timestamp 0
transform 1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_107
timestamp 0
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_138
timestamp 0
transform 1 0 13800 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_150
timestamp 0
transform 1 0 14904 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_162
timestamp 0
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_185
timestamp 0
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_274
timestamp 0
transform 1 0 26312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_57
timestamp 0
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_93
timestamp 0
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_98
timestamp 0
transform 1 0 10120 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_110
timestamp 0
transform 1 0 11224 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_122
timestamp 0
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_134
timestamp 0
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_149
timestamp 0
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_167
timestamp 0
transform 1 0 16468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_179
timestamp 0
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_237
timestamp 0
transform 1 0 22908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 0
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_269
timestamp 0
transform 1 0 25852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 0
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_37
timestamp 0
transform 1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 0
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_65
timestamp 0
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_84
timestamp 0
transform 1 0 8832 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_92
timestamp 0
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_102
timestamp 0
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 0
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_141
timestamp 0
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_178
timestamp 0
transform 1 0 17480 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_186
timestamp 0
transform 1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_220
timestamp 0
transform 1 0 21344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_247
timestamp 0
transform 1 0 23828 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_255
timestamp 0
transform 1 0 24564 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_263
timestamp 0
transform 1 0 25300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_271
timestamp 0
transform 1 0 26036 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 0
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_181
timestamp 0
transform 1 0 17756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 0
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_247
timestamp 0
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 0
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_68
timestamp 0
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_80
timestamp 0
transform 1 0 8464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 0
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_160
timestamp 0
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_173
timestamp 0
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_183
timestamp 0
transform 1 0 17940 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_220
timestamp 0
transform 1 0 21344 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_237
timestamp 0
transform 1 0 22908 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_246
timestamp 0
transform 1 0 23736 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_258
timestamp 0
transform 1 0 24840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_270
timestamp 0
transform 1 0 25944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_276
timestamp 0
transform 1 0 26496 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_23
timestamp 0
transform 1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_51
timestamp 0
transform 1 0 5796 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_68
timestamp 0
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 0
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_113
timestamp 0
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_125
timestamp 0
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 0
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_152
timestamp 0
transform 1 0 15088 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_164
timestamp 0
transform 1 0 16192 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_188
timestamp 0
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_224
timestamp 0
transform 1 0 21712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_232
timestamp 0
transform 1 0 22448 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_236
timestamp 0
transform 1 0 22816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_270
timestamp 0
transform 1 0 25944 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_276
timestamp 0
transform 1 0 26496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_25
timestamp 0
transform 1 0 3404 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_82
timestamp 0
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_148
timestamp 0
transform 1 0 14720 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 0
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_173
timestamp 0
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 0
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 0
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_217
timestamp 0
transform 1 0 21068 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_228
timestamp 0
transform 1 0 22080 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_234
timestamp 0
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_242
timestamp 0
transform 1 0 23368 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_269
timestamp 0
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_7
timestamp 0
transform 1 0 1748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_69
timestamp 0
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_73
timestamp 0
transform 1 0 7820 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_105
timestamp 0
transform 1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_113
timestamp 0
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 0
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_148
timestamp 0
transform 1 0 14720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_179
timestamp 0
transform 1 0 17572 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 0
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_244
timestamp 0
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_253
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_257
timestamp 0
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_266
timestamp 0
transform 1 0 25576 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_11
timestamp 0
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_23
timestamp 0
transform 1 0 3220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_36
timestamp 0
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_40
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 0
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_68
timestamp 0
transform 1 0 7360 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_86
timestamp 0
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_90
timestamp 0
transform 1 0 9384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_148
timestamp 0
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 0
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_201
timestamp 0
transform 1 0 19596 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 0
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_249
timestamp 0
transform 1 0 24012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_257
timestamp 0
transform 1 0 24748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_267
timestamp 0
transform 1 0 25668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_275
timestamp 0
transform 1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_14
timestamp 0
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 0
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_76
timestamp 0
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_93
timestamp 0
transform 1 0 9660 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_105
timestamp 0
transform 1 0 10764 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_117
timestamp 0
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 0
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_183
timestamp 0
transform 1 0 17940 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_213
timestamp 0
transform 1 0 20700 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_226
timestamp 0
transform 1 0 21896 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_238
timestamp 0
transform 1 0 23000 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 0
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_273
timestamp 0
transform 1 0 26220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_30
timestamp 0
transform 1 0 3864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_41
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_47
timestamp 0
transform 1 0 5428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 0
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_60
timestamp 0
transform 1 0 6624 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_72
timestamp 0
transform 1 0 7728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_84
timestamp 0
transform 1 0 8832 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 0
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_144
timestamp 0
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_156
timestamp 0
transform 1 0 15456 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_193
timestamp 0
transform 1 0 18860 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_201
timestamp 0
transform 1 0 19596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_236
timestamp 0
transform 1 0 22816 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_268
timestamp 0
transform 1 0 25760 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_276
timestamp 0
transform 1 0 26496 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 0
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_24
timestamp 0
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_49
timestamp 0
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_69
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_111
timestamp 0
transform 1 0 11316 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_123
timestamp 0
transform 1 0 12420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_129
timestamp 0
transform 1 0 12972 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 0
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_189
timestamp 0
transform 1 0 18492 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 0
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_209
timestamp 0
transform 1 0 20332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_238
timestamp 0
transform 1 0 23000 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 0
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_262
timestamp 0
transform 1 0 25208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_269
timestamp 0
transform 1 0 25852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_11
timestamp 0
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_122
timestamp 0
transform 1 0 12328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_141
timestamp 0
transform 1 0 14076 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_153
timestamp 0
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 0
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_206
timestamp 0
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 0
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_228
timestamp 0
transform 1 0 22080 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_240
timestamp 0
transform 1 0 23184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_252
timestamp 0
transform 1 0 24288 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_275
timestamp 0
transform 1 0 26404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_13
timestamp 0
transform 1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_21
timestamp 0
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_46
timestamp 0
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_58
timestamp 0
transform 1 0 6440 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_68
timestamp 0
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_80
timestamp 0
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_96
timestamp 0
transform 1 0 9936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_110
timestamp 0
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_128
timestamp 0
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_157
timestamp 0
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_162
timestamp 0
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_166
timestamp 0
transform 1 0 16376 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_213
timestamp 0
transform 1 0 20700 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_225
timestamp 0
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_240
timestamp 0
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_253
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_108
timestamp 0
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_123
timestamp 0
transform 1 0 12420 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_131
timestamp 0
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_187
timestamp 0
transform 1 0 18308 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_213
timestamp 0
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 0
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_247
timestamp 0
transform 1 0 23828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_273
timestamp 0
transform 1 0 26220 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 0
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_95
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_107
timestamp 0
transform 1 0 10948 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_119
timestamp 0
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_131
timestamp 0
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_162
timestamp 0
transform 1 0 16008 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_171
timestamp 0
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_183
timestamp 0
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_201
timestamp 0
transform 1 0 19596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_213
timestamp 0
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_217
timestamp 0
transform 1 0 21068 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_241
timestamp 0
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 0
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_14
timestamp 0
transform 1 0 2392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_18
timestamp 0
transform 1 0 2760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_44
timestamp 0
transform 1 0 5152 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_66
timestamp 0
transform 1 0 7176 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_103
timestamp 0
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 0
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_193
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_206
timestamp 0
transform 1 0 20056 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_218
timestamp 0
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_245
timestamp 0
transform 1 0 23644 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_257
timestamp 0
transform 1 0 24748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_263
timestamp 0
transform 1 0 25300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_267
timestamp 0
transform 1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_11
timestamp 0
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_45
timestamp 0
transform 1 0 5244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_80
timestamp 0
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_108
timestamp 0
transform 1 0 11040 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_116
timestamp 0
transform 1 0 11776 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_158
timestamp 0
transform 1 0 15640 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_170
timestamp 0
transform 1 0 16744 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_182
timestamp 0
transform 1 0 17848 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_214
timestamp 0
transform 1 0 20792 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_220
timestamp 0
transform 1 0 21344 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_230
timestamp 0
transform 1 0 22264 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_239
timestamp 0
transform 1 0 23092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_276
timestamp 0
transform 1 0 26496 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_32
timestamp 0
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_44
timestamp 0
transform 1 0 5152 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_80
timestamp 0
transform 1 0 8464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_98
timestamp 0
transform 1 0 10120 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_108
timestamp 0
transform 1 0 11040 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_140
timestamp 0
transform 1 0 13984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 0
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_177
timestamp 0
transform 1 0 17388 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_206
timestamp 0
transform 1 0 20056 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_214
timestamp 0
transform 1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_239
timestamp 0
transform 1 0 23092 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_251
timestamp 0
transform 1 0 24196 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_263
timestamp 0
transform 1 0 25300 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_11
timestamp 0
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_33
timestamp 0
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_42
timestamp 0
transform 1 0 4968 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_54
timestamp 0
transform 1 0 6072 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_72
timestamp 0
transform 1 0 7728 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_179
timestamp 0
transform 1 0 17572 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_212
timestamp 0
transform 1 0 20608 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_244
timestamp 0
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 0
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_31
timestamp 0
transform 1 0 3956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_37
timestamp 0
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_49
timestamp 0
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_103
timestamp 0
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 0
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_136
timestamp 0
transform 1 0 13616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_142
timestamp 0
transform 1 0 14168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 0
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_177
timestamp 0
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_213
timestamp 0
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_245
timestamp 0
transform 1 0 23644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_253
timestamp 0
transform 1 0 24380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_275
timestamp 0
transform 1 0 26404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_20
timestamp 0
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_47
timestamp 0
transform 1 0 5428 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_59
timestamp 0
transform 1 0 6532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_76
timestamp 0
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_89
timestamp 0
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_99
timestamp 0
transform 1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_108
timestamp 0
transform 1 0 11040 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_116
timestamp 0
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_127
timestamp 0
transform 1 0 12788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_168
timestamp 0
transform 1 0 16560 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_180
timestamp 0
transform 1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 0
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_200
timestamp 0
transform 1 0 19504 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_212
timestamp 0
transform 1 0 20608 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_220
timestamp 0
transform 1 0 21344 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_276
timestamp 0
transform 1 0 26496 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_50
timestamp 0
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_83
timestamp 0
transform 1 0 8740 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_155
timestamp 0
transform 1 0 15364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_180
timestamp 0
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_195
timestamp 0
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_207
timestamp 0
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_219
timestamp 0
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 0
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_275
timestamp 0
transform 1 0 26404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_14
timestamp 0
transform 1 0 2392 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_22
timestamp 0
transform 1 0 3128 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_48
timestamp 0
transform 1 0 5520 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_60
timestamp 0
transform 1 0 6624 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 0
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_92
timestamp 0
transform 1 0 9568 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_113
timestamp 0
transform 1 0 11500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_147
timestamp 0
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_164
timestamp 0
transform 1 0 16192 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 0
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_203
timestamp 0
transform 1 0 19780 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_215
timestamp 0
transform 1 0 20884 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_227
timestamp 0
transform 1 0 21988 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_231
timestamp 0
transform 1 0 22356 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_243
timestamp 0
transform 1 0 23460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 0
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_253
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_276
timestamp 0
transform 1 0 26496 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_11
timestamp 0
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_17
timestamp 0
transform 1 0 2668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_27
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_35
timestamp 0
transform 1 0 4324 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_48
timestamp 0
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_60
timestamp 0
transform 1 0 6624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_78
timestamp 0
transform 1 0 8280 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_82
timestamp 0
transform 1 0 8648 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_151
timestamp 0
transform 1 0 14996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_159
timestamp 0
transform 1 0 15732 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_182
timestamp 0
transform 1 0 17848 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_186
timestamp 0
transform 1 0 18216 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_206
timestamp 0
transform 1 0 20056 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_213
timestamp 0
transform 1 0 20700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_221
timestamp 0
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_245
timestamp 0
transform 1 0 23644 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_257
timestamp 0
transform 1 0 24748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_269
timestamp 0
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_25
timestamp 0
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_36
timestamp 0
transform 1 0 4416 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_150
timestamp 0
transform 1 0 14904 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_162
timestamp 0
transform 1 0 16008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_210
timestamp 0
transform 1 0 20424 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_238
timestamp 0
transform 1 0 23000 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_246
timestamp 0
transform 1 0 23736 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_266
timestamp 0
transform 1 0 25576 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_274
timestamp 0
transform 1 0 26312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_11
timestamp 0
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_17
timestamp 0
transform 1 0 2668 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_28
timestamp 0
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_36
timestamp 0
transform 1 0 4416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_40
timestamp 0
transform 1 0 4784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_50
timestamp 0
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_73
timestamp 0
transform 1 0 7820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_85
timestamp 0
transform 1 0 8924 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_100
timestamp 0
transform 1 0 10304 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_129
timestamp 0
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_136
timestamp 0
transform 1 0 13616 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_146
timestamp 0
transform 1 0 14536 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_158
timestamp 0
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 0
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 0
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_228
timestamp 0
transform 1 0 22080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_235
timestamp 0
transform 1 0 22724 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_243
timestamp 0
transform 1 0 23460 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_272
timestamp 0
transform 1 0 26128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_276
timestamp 0
transform 1 0 26496 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_25
timestamp 0
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_38
timestamp 0
transform 1 0 4600 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_42
timestamp 0
transform 1 0 4968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_54
timestamp 0
transform 1 0 6072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_74
timestamp 0
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 0
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_98
timestamp 0
transform 1 0 10120 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_110
timestamp 0
transform 1 0 11224 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_122
timestamp 0
transform 1 0 12328 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_134
timestamp 0
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_145
timestamp 0
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_149
timestamp 0
transform 1 0 14812 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_161
timestamp 0
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_188
timestamp 0
transform 1 0 18400 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_231
timestamp 0
transform 1 0 22356 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_243
timestamp 0
transform 1 0 23460 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_9
timestamp 0
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_26
timestamp 0
transform 1 0 3496 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_65
timestamp 0
transform 1 0 7084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_77
timestamp 0
transform 1 0 8188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_85
timestamp 0
transform 1 0 8924 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_96
timestamp 0
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_108
timestamp 0
transform 1 0 11040 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_122
timestamp 0
transform 1 0 12328 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_134
timestamp 0
transform 1 0 13432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_228
timestamp 0
transform 1 0 22080 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_240
timestamp 0
transform 1 0 23184 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_258
timestamp 0
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_262
timestamp 0
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_269
timestamp 0
transform 1 0 25852 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_18
timestamp 0
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 0
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_37
timestamp 0
transform 1 0 4508 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_42
timestamp 0
transform 1 0 4968 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_49
timestamp 0
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_61
timestamp 0
transform 1 0 6716 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_75
timestamp 0
transform 1 0 8004 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_101
timestamp 0
transform 1 0 10396 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_107
timestamp 0
transform 1 0 10948 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_124
timestamp 0
transform 1 0 12512 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_136
timestamp 0
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_160
timestamp 0
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_230
timestamp 0
transform 1 0 22264 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_238
timestamp 0
transform 1 0 23000 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_256
timestamp 0
transform 1 0 24656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_268
timestamp 0
transform 1 0 25760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_276
timestamp 0
transform 1 0 26496 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_11
timestamp 0
transform 1 0 2116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_16
timestamp 0
transform 1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_34
timestamp 0
transform 1 0 4232 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_46
timestamp 0
transform 1 0 5336 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 0
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_83
timestamp 0
transform 1 0 8740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_142
timestamp 0
transform 1 0 14168 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_156
timestamp 0
transform 1 0 15456 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_175
timestamp 0
transform 1 0 17204 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_221
timestamp 0
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_236
timestamp 0
transform 1 0 22816 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_244
timestamp 0
transform 1 0 23552 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_265
timestamp 0
transform 1 0 25484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_273
timestamp 0
transform 1 0 26220 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_25
timestamp 0
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_37
timestamp 0
transform 1 0 4508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_63
timestamp 0
transform 1 0 6900 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_93
timestamp 0
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_157
timestamp 0
transform 1 0 15548 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_219
timestamp 0
transform 1 0 21252 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_227
timestamp 0
transform 1 0 21988 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_259
timestamp 0
transform 1 0 24932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_271
timestamp 0
transform 1 0 26036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_66
timestamp 0
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_79
timestamp 0
transform 1 0 8372 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_91
timestamp 0
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_103
timestamp 0
transform 1 0 10580 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_153
timestamp 0
transform 1 0 15180 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_210
timestamp 0
transform 1 0 20424 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 0
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_229
timestamp 0
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_263
timestamp 0
transform 1 0 25300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_275
timestamp 0
transform 1 0 26404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_7
timestamp 0
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_24
timestamp 0
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_37
timestamp 0
transform 1 0 4508 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_57
timestamp 0
transform 1 0 6348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_69
timestamp 0
transform 1 0 7452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 0
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 0
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_121
timestamp 0
transform 1 0 12236 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_129
timestamp 0
transform 1 0 12972 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_134
timestamp 0
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 0
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 0
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 0
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 0
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_203
timestamp 0
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_230
timestamp 0
transform 1 0 22264 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_238
timestamp 0
transform 1 0 23000 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 0
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_256
timestamp 0
transform 1 0 24656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_268
timestamp 0
transform 1 0 25760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_276
timestamp 0
transform 1 0 26496 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_11
timestamp 0
transform 1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_16
timestamp 0
transform 1 0 2576 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_26
timestamp 0
transform 1 0 3496 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_38
timestamp 0
transform 1 0 4600 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_44
timestamp 0
transform 1 0 5152 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_48
timestamp 0
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_66
timestamp 0
transform 1 0 7176 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_78
timestamp 0
transform 1 0 8280 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_89
timestamp 0
transform 1 0 9292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_97
timestamp 0
transform 1 0 10028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_107
timestamp 0
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 0
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 0
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 0
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 0
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 0
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_193
timestamp 0
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_208
timestamp 0
transform 1 0 20240 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_220
timestamp 0
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 0
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 0
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 0
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_273
timestamp 0
transform 1 0 26220 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 0
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_41
timestamp 0
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_45
timestamp 0
transform 1 0 5244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_62
timestamp 0
transform 1 0 6808 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_88
timestamp 0
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_98
timestamp 0
transform 1 0 10120 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_122
timestamp 0
transform 1 0 12328 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_128
timestamp 0
transform 1 0 12880 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 0
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_153
timestamp 0
transform 1 0 15180 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_166
timestamp 0
transform 1 0 16376 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_174
timestamp 0
transform 1 0 17112 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_178
timestamp 0
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_190
timestamp 0
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_204
timestamp 0
transform 1 0 19872 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_218
timestamp 0
transform 1 0 21160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_229
timestamp 0
transform 1 0 22172 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_235
timestamp 0
transform 1 0 22724 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_242
timestamp 0
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 0
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_63
timestamp 0
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_80
timestamp 0
transform 1 0 8464 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_116
timestamp 0
transform 1 0 11776 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_128
timestamp 0
transform 1 0 12880 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_149
timestamp 0
transform 1 0 14812 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 0
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_185
timestamp 0
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_189
timestamp 0
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_202
timestamp 0
transform 1 0 19688 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_228
timestamp 0
transform 1 0 22080 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_252
timestamp 0
transform 1 0 24288 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_264
timestamp 0
transform 1 0 25392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_276
timestamp 0
transform 1 0 26496 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_33
timestamp 0
transform 1 0 4140 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_52
timestamp 0
transform 1 0 5888 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_64
timestamp 0
transform 1 0 6992 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_94
timestamp 0
transform 1 0 9752 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_121
timestamp 0
transform 1 0 12236 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 0
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 0
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_220
timestamp 0
transform 1 0 21344 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_232
timestamp 0
transform 1 0 22448 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_243
timestamp 0
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 0
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 0
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_43
timestamp 0
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_83
timestamp 0
transform 1 0 8740 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 0
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_130
timestamp 0
transform 1 0 13064 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_149
timestamp 0
transform 1 0 14812 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_153
timestamp 0
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_186
timestamp 0
transform 1 0 18216 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_211
timestamp 0
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 0
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 0
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 0
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_273
timestamp 0
transform 1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 0
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 0
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_57
timestamp 0
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_69
timestamp 0
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 0
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_93
timestamp 0
transform 1 0 9660 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_97
timestamp 0
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_104
timestamp 0
transform 1 0 10672 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_111
timestamp 0
transform 1 0 11316 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_113
timestamp 0
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_118
timestamp 0
transform 1 0 11960 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_125
timestamp 0
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 0
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_146
timestamp 0
transform 1 0 14536 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_158
timestamp 0
transform 1 0 15640 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_166
timestamp 0
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_169
timestamp 0
transform 1 0 16652 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_177
timestamp 0
transform 1 0 17388 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 0
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 0
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_203
timestamp 0
transform 1 0 19780 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_209
timestamp 0
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 0
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 0
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 0
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 0
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 17388 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 7084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform 1 0 12236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform 1 0 20700 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 0
transform -1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 0
transform -1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 0
transform 1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 0
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 0
transform -1 0 16560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 0
transform 1 0 12972 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform -1 0 26588 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output11
timestamp 0
transform -1 0 20332 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output12
timestamp 0
transform -1 0 11316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output13
timestamp 0
transform -1 0 10672 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output14
timestamp 0
transform -1 0 10028 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output15
timestamp 0
transform -1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output16
timestamp 0
transform -1 0 12604 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output17
timestamp 0
transform -1 0 17756 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output18
timestamp 0
transform -1 0 14536 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output19
timestamp 0
transform 1 0 26312 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output20
timestamp 0
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_47
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 26864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_48
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 26864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_49
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 26864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_50
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 26864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_51
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_52
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 26864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_53
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_54
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 26864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_55
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_56
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 26864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_57
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_58
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 26864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_59
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 26864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_60
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 26864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_61
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 26864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_62
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 26864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_63
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 26864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_64
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 26864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_65
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 26864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_66
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 26864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_67
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 26864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_68
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 26864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_69
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 26864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_70
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 26864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_71
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 26864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_72
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 26864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_73
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 26864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_74
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 26864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_75
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 26864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_76
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 26864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_77
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 26864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_78
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 26864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_79
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 26864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_80
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 26864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_81
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 26864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_82
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 26864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_83
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 26864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_84
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 26864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_85
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 26864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_86
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 0
transform -1 0 26864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_87
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 0
transform -1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_88
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 0
transform -1 0 26864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_89
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 0
transform -1 0 26864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_90
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 0
transform -1 0 26864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_91
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 0
transform -1 0 26864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_92
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 0
transform -1 0 26864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_93
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 0
transform -1 0 26864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_94
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_95
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_97
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_103
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_104
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_105
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_106
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_107
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_108
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_109
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_110
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_111
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_112
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_113
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_114
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_115
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_116
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_117
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_118
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_119
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_120
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_121
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_122
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_123
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_124
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_125
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_126
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_127
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_128
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_129
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_130
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_131
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_132
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_133
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_134
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_135
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_136
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_137
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_138
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_139
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_140
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_141
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_142
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_144
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_145
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_146
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_147
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_149
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_150
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_151
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_155
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_156
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_160
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_170
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_175
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_176
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_179
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_180
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_181
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_184
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_185
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_186
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_187
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_189
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_190
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_191
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_192
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_194
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_195
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_196
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_200
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_201
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_205
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_215
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_220
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_221
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_224
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_225
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_226
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_229
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_230
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_231
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_232
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_233
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_234
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_235
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_236
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_237
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_238
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_239
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_240
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_241
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_242
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_243
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_244
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_245
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_246
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_247
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_248
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_249
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_250
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_251
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_252
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_253
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_254
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_255
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_256
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_257
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_258
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_259
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_260
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_261
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_262
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_263
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_264
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_265
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_266
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_267
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_268
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_269
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_270
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_271
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_272
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_273
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_274
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_275
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_276
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_277
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_278
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_279
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_280
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_281
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_282
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_283
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_284
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_285
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_286
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_287
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_288
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_289
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_290
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_291
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_292
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_293
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_294
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_295
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_296
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_297
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_298
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_299
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_300
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_301
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_302
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_303
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_304
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_305
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_306
timestamp 0
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_307
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_308
timestamp 0
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_309
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_310
timestamp 0
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_311
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_312
timestamp 0
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_313
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
<< labels >>
rlabel metal1 s 13984 27200 13984 27200 4 VGND
rlabel metal1 s 13984 27744 13984 27744 4 VPWR
rlabel metal1 s 21528 16966 21528 16966 4 _0000_
rlabel metal1 s 25813 17238 25813 17238 4 _0001_
rlabel metal1 s 26135 17578 26135 17578 4 _0002_
rlabel metal1 s 23375 17578 23375 17578 4 _0003_
rlabel metal1 s 22908 16218 22908 16218 4 _0004_
rlabel metal2 s 22218 19142 22218 19142 4 _0005_
rlabel metal2 s 26266 18530 26266 18530 4 _0006_
rlabel metal2 s 25714 21080 25714 21080 4 _0007_
rlabel metal1 s 24518 17850 24518 17850 4 _0008_
rlabel metal2 s 23874 18088 23874 18088 4 _0009_
rlabel metal1 s 20332 26758 20332 26758 4 _0010_
rlabel metal1 s 11967 25194 11967 25194 4 _0011_
rlabel metal1 s 11875 26282 11875 26282 4 _0012_
rlabel metal1 s 11454 25738 11454 25738 4 _0013_
rlabel metal1 s 11316 23494 11316 23494 4 _0014_
rlabel metal1 s 12151 23018 12151 23018 4 _0015_
rlabel metal1 s 16468 26758 16468 26758 4 _0016_
rlabel metal2 s 14674 26350 14674 26350 4 _0017_
rlabel metal1 s 17756 22678 17756 22678 4 _0018_
rlabel metal2 s 18998 22848 18998 22848 4 _0019_
rlabel metal1 s 21903 24106 21903 24106 4 _0020_
rlabel metal1 s 21443 25942 21443 25942 4 _0021_
rlabel metal2 s 21942 10166 21942 10166 4 _0022_
rlabel metal1 s 25951 15402 25951 15402 4 _0023_
rlabel metal2 s 22862 15198 22862 15198 4 _0024_
rlabel metal2 s 26358 14654 26358 14654 4 _0025_
rlabel metal1 s 22915 14314 22915 14314 4 _0026_
rlabel metal1 s 23191 9962 23191 9962 4 _0027_
rlabel metal1 s 26227 13294 26227 13294 4 _0028_
rlabel metal2 s 25162 14552 25162 14552 4 _0029_
rlabel metal1 s 24610 13974 24610 13974 4 _0030_
rlabel metal1 s 22954 13498 22954 13498 4 _0031_
rlabel metal1 s 21765 19754 21765 19754 4 _0032_
rlabel metal2 s 24518 22814 24518 22814 4 _0033_
rlabel metal1 s 24387 23018 24387 23018 4 _0034_
rlabel metal2 s 24518 23902 24518 23902 4 _0035_
rlabel metal1 s 23414 26282 23414 26282 4 _0036_
rlabel metal2 s 25806 8296 25806 8296 4 _0037_
rlabel metal2 s 24518 3196 24518 3196 4 _0038_
rlabel metal2 s 24978 3944 24978 3944 4 _0039_
rlabel metal2 s 22586 4318 22586 4318 4 _0040_
rlabel metal2 s 21758 11560 21758 11560 4 _0041_
rlabel metal2 s 25714 11288 25714 11288 4 _0042_
rlabel metal1 s 25123 11798 25123 11798 4 _0043_
rlabel metal1 s 22639 12138 22639 12138 4 _0044_
rlabel metal1 s 22540 3162 22540 3162 4 _0045_
rlabel metal1 s 19688 25466 19688 25466 4 _0046_
rlabel metal1 s 10718 24922 10718 24922 4 _0047_
rlabel metal1 s 10488 26282 10488 26282 4 _0048_
rlabel metal1 s 11132 25942 11132 25942 4 _0049_
rlabel metal1 s 10120 22542 10120 22542 4 _0050_
rlabel metal1 s 11132 22746 11132 22746 4 _0051_
rlabel metal2 s 18078 26112 18078 26112 4 _0052_
rlabel metal1 s 13340 25942 13340 25942 4 _0053_
rlabel metal1 s 16514 23596 16514 23596 4 _0054_
rlabel metal2 s 19458 22814 19458 22814 4 _0055_
rlabel metal1 s 20240 24106 20240 24106 4 _0056_
rlabel metal1 s 20792 24718 20792 24718 4 _0057_
rlabel metal2 s 22034 20060 22034 20060 4 _0058_
rlabel metal1 s 24012 22202 24012 22202 4 _0059_
rlabel metal1 s 22770 22984 22770 22984 4 _0060_
rlabel metal1 s 23598 23766 23598 23766 4 _0061_
rlabel metal1 s 22310 25398 22310 25398 4 _0062_
rlabel metal2 s 24702 7548 24702 7548 4 _0063_
rlabel metal1 s 23460 3094 23460 3094 4 _0064_
rlabel metal1 s 24380 4182 24380 4182 4 _0065_
rlabel metal2 s 22126 4318 22126 4318 4 _0066_
rlabel metal2 s 20194 11934 20194 11934 4 _0067_
rlabel metal2 s 24702 10914 24702 10914 4 _0068_
rlabel metal1 s 23644 11798 23644 11798 4 _0069_
rlabel metal1 s 21528 12614 21528 12614 4 _0070_
rlabel metal1 s 21574 3570 21574 3570 4 _0071_
rlabel metal1 s 18722 26010 18722 26010 4 _0072_
rlabel metal1 s 8321 25194 8321 25194 4 _0073_
rlabel metal2 s 7130 26078 7130 26078 4 _0074_
rlabel metal2 s 7677 26350 7677 26350 4 _0075_
rlabel metal1 s 8786 21896 8786 21896 4 _0076_
rlabel metal2 s 11178 21794 11178 21794 4 _0077_
rlabel metal1 s 17710 25466 17710 25466 4 _0078_
rlabel metal2 s 12737 26350 12737 26350 4 _0079_
rlabel metal1 s 14117 13974 14117 13974 4 _0080_
rlabel metal2 s 2346 22882 2346 22882 4 _0081_
rlabel metal2 s 2341 21522 2341 21522 4 _0082_
rlabel metal1 s 6739 22746 6739 22746 4 _0083_
rlabel metal1 s 1610 6664 1610 6664 4 _0084_
rlabel metal1 s 9000 19754 9000 19754 4 _0085_
rlabel metal1 s 16049 5270 16049 5270 4 _0086_
rlabel metal1 s 12088 10642 12088 10642 4 _0087_
rlabel metal1 s 20056 15130 20056 15130 4 _0088_
rlabel metal1 s 6516 12886 6516 12886 4 _0089_
rlabel metal2 s 8146 15470 8146 15470 4 _0090_
rlabel metal2 s 2893 4182 2893 4182 4 _0091_
rlabel metal2 s 1886 6494 1886 6494 4 _0092_
rlabel metal1 s 6568 16082 6568 16082 4 _0093_
rlabel metal1 s 19197 10710 19197 10710 4 _0094_
rlabel metal1 s 12047 9962 12047 9962 4 _0095_
rlabel metal1 s 20056 12954 20056 12954 4 _0096_
rlabel metal2 s 4646 12002 4646 12002 4 _0097_
rlabel metal2 s 4738 21726 4738 21726 4 _0098_
rlabel metal1 s 4457 4182 4457 4182 4 _0099_
rlabel metal1 s 7263 7854 7263 7854 4 _0100_
rlabel metal2 s 6762 20706 6762 20706 4 _0101_
rlabel metal1 s 14536 21114 14536 21114 4 _0102_
rlabel metal1 s 13836 5202 13836 5202 4 _0103_
rlabel metal1 s 14520 16150 14520 16150 4 _0104_
rlabel metal1 s 2244 23698 2244 23698 4 _0105_
rlabel metal1 s 5239 24106 5239 24106 4 _0106_
rlabel metal2 s 4641 23766 4641 23766 4 _0107_
rlabel metal1 s 9138 8534 9138 8534 4 _0108_
rlabel metal2 s 6578 19618 6578 19618 4 _0109_
rlabel metal2 s 14398 22882 14398 22882 4 _0110_
rlabel metal2 s 12093 7446 12093 7446 4 _0111_
rlabel metal1 s 17940 16218 17940 16218 4 _0112_
rlabel metal2 s 2157 24174 2157 24174 4 _0113_
rlabel metal1 s 3726 26214 3726 26214 4 _0114_
rlabel metal1 s 4779 26282 4779 26282 4 _0115_
rlabel metal2 s 2162 11526 2162 11526 4 _0116_
rlabel metal1 s 9598 18666 9598 18666 4 _0117_
rlabel metal1 s 14669 26282 14669 26282 4 _0118_
rlabel metal1 s 13002 23766 13002 23766 4 _0119_
rlabel metal1 s 14290 13226 14290 13226 4 _0120_
rlabel metal1 s 1973 17646 1973 17646 4 _0121_
rlabel metal2 s 2254 16966 2254 16966 4 _0122_
rlabel metal1 s 7999 10642 7999 10642 4 _0123_
rlabel metal1 s 1789 8942 1789 8942 4 _0124_
rlabel metal1 s 6660 18258 6660 18258 4 _0125_
rlabel metal2 s 15221 10710 15221 10710 4 _0126_
rlabel metal1 s 13013 12886 13013 12886 4 _0127_
rlabel metal1 s 19876 13226 19876 13226 4 _0128_
rlabel metal2 s 2801 18258 2801 18258 4 _0129_
rlabel metal2 s 3358 15674 3358 15674 4 _0130_
rlabel metal1 s 6716 5882 6716 5882 4 _0131_
rlabel metal1 s 3951 9554 3951 9554 4 _0132_
rlabel metal2 s 11546 19618 11546 19618 4 _0133_
rlabel metal2 s 18818 9962 18818 9962 4 _0134_
rlabel metal1 s 13105 19822 13105 19822 4 _0135_
rlabel metal1 s 14490 16218 14490 16218 4 _0136_
rlabel metal2 s 2438 19618 2438 19618 4 _0137_
rlabel metal2 s 2438 20706 2438 20706 4 _0138_
rlabel metal2 s 6757 6766 6757 6766 4 _0139_
rlabel metal1 s 1876 5678 1876 5678 4 _0140_
rlabel metal1 s 11720 16082 11720 16082 4 _0141_
rlabel metal1 s 14888 7446 14888 7446 4 _0142_
rlabel metal1 s 13059 19414 13059 19414 4 _0143_
rlabel metal2 s 15134 18530 15134 18530 4 _0144_
rlabel metal2 s 12558 13498 12558 13498 4 _0145_
rlabel metal1 s 5791 25262 5791 25262 4 _0146_
rlabel metal1 s 8433 23018 8433 23018 4 _0147_
rlabel metal1 s 6297 8874 6297 8874 4 _0148_
rlabel metal2 s 6941 17646 6941 17646 4 _0149_
rlabel metal1 s 15364 25466 15364 25466 4 _0150_
rlabel metal1 s 13013 23086 13013 23086 4 _0151_
rlabel metal2 s 15778 13702 15778 13702 4 _0152_
rlabel metal2 s 2157 12138 2157 12138 4 _0153_
rlabel metal1 s 3312 14586 3312 14586 4 _0154_
rlabel metal2 s 7222 3298 7222 3298 4 _0155_
rlabel metal2 s 2714 9350 2714 9350 4 _0156_
rlabel metal1 s 4411 3026 4411 3026 4 _0157_
rlabel metal2 s 15318 9826 15318 9826 4 _0158_
rlabel metal1 s 12231 3026 12231 3026 4 _0159_
rlabel metal1 s 17878 17238 17878 17238 4 _0160_
rlabel metal1 s 8684 12818 8684 12818 4 _0161_
rlabel metal1 s 4871 18326 4871 18326 4 _0162_
rlabel metal1 s 7028 4114 7028 4114 4 _0163_
rlabel metal1 s 3986 6698 3986 6698 4 _0164_
rlabel metal1 s 11898 16490 11898 16490 4 _0165_
rlabel metal1 s 15451 6766 15451 6766 4 _0166_
rlabel metal1 s 11868 5882 11868 5882 4 _0167_
rlabel metal1 s 16866 12886 16866 12886 4 _0168_
rlabel metal2 s 2806 13022 2806 13022 4 _0169_
rlabel metal2 s 2162 15606 2162 15606 4 _0170_
rlabel metal1 s 9420 3502 9420 3502 4 _0171_
rlabel metal1 s 3848 8874 3848 8874 4 _0172_
rlabel metal2 s 5934 15266 5934 15266 4 _0173_
rlabel metal2 s 15410 3298 15410 3298 4 _0174_
rlabel metal1 s 12921 4522 12921 4522 4 _0175_
rlabel metal1 s 15778 16218 15778 16218 4 _0176_
rlabel metal2 s 9430 12002 9430 12002 4 _0177_
rlabel metal1 s 9138 15402 9138 15402 4 _0178_
rlabel metal2 s 10630 4114 10630 4114 4 _0179_
rlabel metal1 s 9506 7786 9506 7786 4 _0180_
rlabel metal1 s 10161 16558 10161 16558 4 _0181_
rlabel metal1 s 18507 3094 18507 3094 4 _0182_
rlabel metal1 s 13478 8058 13478 8058 4 _0183_
rlabel metal1 s 17004 13226 17004 13226 4 _0184_
rlabel metal2 s 6394 12002 6394 12002 4 _0185_
rlabel metal2 s 8781 14994 8781 14994 4 _0186_
rlabel metal1 s 9322 3094 9322 3094 4 _0187_
rlabel metal1 s 6568 9554 6568 9554 4 _0188_
rlabel metal1 s 5561 3434 5561 3434 4 _0189_
rlabel metal2 s 16330 3298 16330 3298 4 _0190_
rlabel metal2 s 12461 3502 12461 3502 4 _0191_
rlabel metal1 s 19922 17238 19922 17238 4 _0192_
rlabel metal2 s 11090 12818 11090 12818 4 _0193_
rlabel metal2 s 9287 18326 9287 18326 4 _0194_
rlabel metal2 s 9793 6290 9793 6290 4 _0195_
rlabel metal1 s 9414 9962 9414 9962 4 _0196_
rlabel metal1 s 11766 15470 11766 15470 4 _0197_
rlabel metal1 s 18266 8942 18266 8942 4 _0198_
rlabel metal1 s 12174 7786 12174 7786 4 _0199_
rlabel metal1 s 22402 8942 22402 8942 4 _0200_
rlabel metal1 s 22724 7922 22724 7922 4 _0201_
rlabel metal1 s 23874 8840 23874 8840 4 _0202_
rlabel metal1 s 24886 6766 24886 6766 4 _0203_
rlabel metal1 s 25024 8874 25024 8874 4 _0204_
rlabel metal1 s 24012 9146 24012 9146 4 _0205_
rlabel metal2 s 19826 8126 19826 8126 4 _0206_
rlabel metal1 s 25024 6086 25024 6086 4 _0207_
rlabel metal1 s 25668 9554 25668 9554 4 _0208_
rlabel metal2 s 25622 5950 25622 5950 4 _0209_
rlabel metal2 s 25254 8262 25254 8262 4 _0210_
rlabel metal2 s 25806 10812 25806 10812 4 _0211_
rlabel metal1 s 25346 8976 25346 8976 4 _0212_
rlabel metal2 s 24978 9520 24978 9520 4 _0213_
rlabel metal2 s 23966 9146 23966 9146 4 _0214_
rlabel metal1 s 23782 8398 23782 8398 4 _0215_
rlabel metal1 s 23920 8602 23920 8602 4 _0216_
rlabel metal1 s 23552 8942 23552 8942 4 _0217_
rlabel metal1 s 25438 8908 25438 8908 4 _0218_
rlabel metal1 s 22632 9486 22632 9486 4 _0219_
rlabel metal2 s 25622 9146 25622 9146 4 _0220_
rlabel metal1 s 23828 8534 23828 8534 4 _0221_
rlabel metal1 s 19596 7854 19596 7854 4 _0222_
rlabel metal1 s 20792 5746 20792 5746 4 _0223_
rlabel metal2 s 20654 6562 20654 6562 4 _0224_
rlabel metal2 s 21942 5338 21942 5338 4 _0225_
rlabel metal2 s 21390 11390 21390 11390 4 _0226_
rlabel metal2 s 22034 12342 22034 12342 4 _0227_
rlabel metal1 s 24426 10778 24426 10778 4 _0228_
rlabel metal1 s 24196 12206 24196 12206 4 _0229_
rlabel metal2 s 25162 10404 25162 10404 4 _0230_
rlabel metal1 s 24702 10642 24702 10642 4 _0231_
rlabel metal2 s 21574 9826 21574 9826 4 _0232_
rlabel metal2 s 20838 11764 20838 11764 4 _0233_
rlabel metal2 s 22218 5066 22218 5066 4 _0234_
rlabel metal1 s 25714 5780 25714 5780 4 _0235_
rlabel metal1 s 24932 4590 24932 4590 4 _0236_
rlabel metal1 s 24104 4590 24104 4590 4 _0237_
rlabel metal2 s 25530 20876 25530 20876 4 _0238_
rlabel metal1 s 25254 19754 25254 19754 4 _0239_
rlabel metal2 s 24702 20196 24702 20196 4 _0240_
rlabel metal1 s 23690 19958 23690 19958 4 _0241_
rlabel metal1 s 25254 20332 25254 20332 4 _0242_
rlabel metal1 s 25070 20570 25070 20570 4 _0243_
rlabel metal1 s 24564 20434 24564 20434 4 _0244_
rlabel metal1 s 24646 20298 24646 20298 4 _0245_
rlabel metal1 s 24288 20910 24288 20910 4 _0246_
rlabel metal1 s 23828 20026 23828 20026 4 _0247_
rlabel metal2 s 24150 20638 24150 20638 4 _0248_
rlabel metal2 s 21758 21828 21758 21828 4 _0249_
rlabel metal1 s 23460 22134 23460 22134 4 _0250_
rlabel metal1 s 9154 22610 9154 22610 4 _0251_
rlabel metal2 s 19734 18972 19734 18972 4 _0252_
rlabel metal1 s 20654 21556 20654 21556 4 _0253_
rlabel metal1 s 20102 20434 20102 20434 4 _0254_
rlabel metal1 s 20930 19482 20930 19482 4 _0255_
rlabel metal2 s 19366 16167 19366 16167 4 _0256_
rlabel metal2 s 21666 25772 21666 25772 4 _0257_
rlabel metal2 s 20470 20638 20470 20638 4 _0258_
rlabel metal1 s 16836 21998 16836 21998 4 _0259_
rlabel metal2 s 22402 23426 22402 23426 4 _0260_
rlabel metal2 s 22862 23868 22862 23868 4 _0261_
rlabel metal2 s 23230 23868 23230 23868 4 _0262_
rlabel metal1 s 21666 22066 21666 22066 4 _0263_
rlabel metal2 s 22310 22372 22310 22372 4 _0264_
rlabel metal1 s 22494 22746 22494 22746 4 _0265_
rlabel metal1 s 20056 20230 20056 20230 4 _0266_
rlabel metal2 s 23506 21658 23506 21658 4 _0267_
rlabel metal1 s 24104 21862 24104 21862 4 _0268_
rlabel metal2 s 22218 20570 22218 20570 4 _0269_
rlabel metal1 s 21666 20434 21666 20434 4 _0270_
rlabel metal1 s 19734 23290 19734 23290 4 _0271_
rlabel metal2 s 19918 24446 19918 24446 4 _0272_
rlabel metal1 s 20194 23834 20194 23834 4 _0273_
rlabel metal2 s 19458 23290 19458 23290 4 _0274_
rlabel metal1 s 10258 23086 10258 23086 4 _0275_
rlabel metal1 s 18078 18768 18078 18768 4 _0276_
rlabel metal2 s 17710 18258 17710 18258 4 _0277_
rlabel metal1 s 20010 16082 20010 16082 4 _0278_
rlabel metal1 s 17250 19380 17250 19380 4 _0279_
rlabel metal1 s 5152 23018 5152 23018 4 _0280_
rlabel metal1 s 13892 9146 13892 9146 4 _0281_
rlabel metal1 s 13662 17170 13662 17170 4 _0282_
rlabel metal1 s 14628 9690 14628 9690 4 _0283_
rlabel metal2 s 17894 19210 17894 19210 4 _0284_
rlabel metal2 s 14490 11084 14490 11084 4 _0285_
rlabel metal2 s 4002 22372 4002 22372 4 _0286_
rlabel metal1 s 18354 15402 18354 15402 4 _0287_
rlabel metal2 s 13754 10336 13754 10336 4 _0288_
rlabel metal3 s 18354 20349 18354 20349 4 _0289_
rlabel metal1 s 18446 13226 18446 13226 4 _0290_
rlabel metal1 s 17066 4624 17066 4624 4 _0291_
rlabel metal1 s 16790 14382 16790 14382 4 _0292_
rlabel metal1 s 14030 4250 14030 4250 4 _0293_
rlabel metal2 s 14766 7684 14766 7684 4 _0294_
rlabel metal1 s 19136 20842 19136 20842 4 _0295_
rlabel metal1 s 15962 17136 15962 17136 4 _0296_
rlabel metal1 s 8464 22678 8464 22678 4 _0297_
rlabel metal1 s 5336 23086 5336 23086 4 _0298_
rlabel metal1 s 13800 20434 13800 20434 4 _0299_
rlabel metal1 s 14214 20230 14214 20230 4 _0300_
rlabel metal2 s 14674 10234 14674 10234 4 _0301_
rlabel metal2 s 12512 19924 12512 19924 4 _0302_
rlabel metal2 s 9154 22304 9154 22304 4 _0303_
rlabel metal1 s 13938 26996 13938 26996 4 _0304_
rlabel metal1 s 17250 8058 17250 8058 4 _0305_
rlabel metal1 s 17388 9690 17388 9690 4 _0306_
rlabel metal1 s 17158 10234 17158 10234 4 _0307_
rlabel metal1 s 15686 22202 15686 22202 4 _0308_
rlabel metal3 s 17342 10659 17342 10659 4 _0309_
rlabel metal1 s 17434 4250 17434 4250 4 _0310_
rlabel metal1 s 16974 4794 16974 4794 4 _0311_
rlabel metal2 s 16974 10234 16974 10234 4 _0312_
rlabel metal3 s 17526 10251 17526 10251 4 _0313_
rlabel metal2 s 17526 26350 17526 26350 4 _0314_
rlabel metal2 s 13846 16932 13846 16932 4 _0315_
rlabel metal2 s 13018 17986 13018 17986 4 _0316_
rlabel metal1 s 10396 17850 10396 17850 4 _0317_
rlabel metal1 s 7636 16422 7636 16422 4 _0318_
rlabel metal1 s 8832 18938 8832 18938 4 _0319_
rlabel metal1 s 6624 19414 6624 19414 4 _0320_
rlabel metal1 s 8694 19278 8694 19278 4 _0321_
rlabel metal1 s 10718 18734 10718 18734 4 _0322_
rlabel metal1 s 11960 22610 11960 22610 4 _0323_
rlabel metal1 s 12144 22610 12144 22610 4 _0324_
rlabel metal2 s 11454 8228 11454 8228 4 _0325_
rlabel metal2 s 10534 9622 10534 9622 4 _0326_
rlabel metal1 s 6256 10030 6256 10030 4 _0327_
rlabel metal2 s 6118 10336 6118 10336 4 _0328_
rlabel metal1 s 4646 10642 4646 10642 4 _0329_
rlabel metal1 s 6026 9996 6026 9996 4 _0330_
rlabel metal2 s 5290 6970 5290 6970 4 _0331_
rlabel metal2 s 5934 6681 5934 6681 4 _0332_
rlabel metal1 s 10718 10574 10718 10574 4 _0333_
rlabel metal1 s 10074 22950 10074 22950 4 _0334_
rlabel metal2 s 9522 22916 9522 22916 4 _0335_
rlabel metal4 s 5405 22100 5405 22100 4 _0336_
rlabel metal2 s 9614 10812 9614 10812 4 _0337_
rlabel metal1 s 9338 4794 9338 4794 4 _0338_
rlabel metal1 s 8786 22406 8786 22406 4 _0339_
rlabel metal2 s 6026 4998 6026 4998 4 _0340_
rlabel metal1 s 8694 5338 8694 5338 4 _0341_
rlabel metal1 s 10672 4454 10672 4454 4 _0342_
rlabel metal1 s 8878 6358 8878 6358 4 _0343_
rlabel metal2 s 9430 8534 9430 8534 4 _0344_
rlabel metal3 s 10557 26860 10557 26860 4 _0345_
rlabel metal1 s 10120 25670 10120 25670 4 _0346_
rlabel metal1 s 10718 15130 10718 15130 4 _0347_
rlabel metal1 s 10258 15606 10258 15606 4 _0348_
rlabel metal2 s 5934 21692 5934 21692 4 _0349_
rlabel metal1 s 6532 22950 6532 22950 4 _0350_
rlabel metal1 s 4462 15674 4462 15674 4 _0351_
rlabel metal1 s 5474 16762 5474 16762 4 _0352_
rlabel metal1 s 5382 20298 5382 20298 4 _0353_
rlabel metal1 s 6210 21624 6210 21624 4 _0354_
rlabel metal1 s 7636 20910 7636 20910 4 _0355_
rlabel metal1 s 10166 21114 10166 21114 4 _0356_
rlabel metal1 s 10028 26962 10028 26962 4 _0357_
rlabel metal1 s 11638 11866 11638 11866 4 _0358_
rlabel metal1 s 10902 13901 10902 13901 4 _0359_
rlabel metal2 s 5934 12580 5934 12580 4 _0360_
rlabel metal1 s 7728 12682 7728 12682 4 _0361_
rlabel metal1 s 4370 22406 4370 22406 4 _0362_
rlabel metal1 s 5750 13396 5750 13396 4 _0363_
rlabel metal2 s 4830 19210 4830 19210 4 _0364_
rlabel metal2 s 5658 14773 5658 14773 4 _0365_
rlabel metal1 s 6762 13430 6762 13430 4 _0366_
rlabel metal2 s 10442 15827 10442 15827 4 _0367_
rlabel metal2 s 10350 24956 10350 24956 4 _0368_
rlabel metal1 s 16330 14348 16330 14348 4 _0369_
rlabel metal1 s 17802 14586 17802 14586 4 _0370_
rlabel metal1 s 20194 16218 20194 16218 4 _0371_
rlabel metal1 s 19550 15674 19550 15674 4 _0372_
rlabel metal1 s 18952 13498 18952 13498 4 _0373_
rlabel metal1 s 18538 14518 18538 14518 4 _0374_
rlabel metal2 s 16698 16524 16698 16524 4 _0375_
rlabel metal2 s 17342 16320 17342 16320 4 _0376_
rlabel metal1 s 18998 16116 18998 16116 4 _0377_
rlabel metal1 s 20010 15946 20010 15946 4 _0378_
rlabel metal1 s 18998 25262 18998 25262 4 _0379_
rlabel metal1 s 22448 24174 22448 24174 4 _0380_
rlabel metal1 s 21873 17170 21873 17170 4 _0381_
rlabel metal1 s 12374 23188 12374 23188 4 _0382_
rlabel metal1 s 21482 9418 21482 9418 4 _0383_
rlabel metal1 s 23644 13294 23644 13294 4 _0384_
rlabel metal2 s 19366 14790 19366 14790 4 _0385_
rlabel metal2 s 21114 5474 21114 5474 4 _0386_
rlabel metal1 s 18791 6834 18791 6834 4 _0387_
rlabel metal1 s 8832 24718 8832 24718 4 _0388_
rlabel metal1 s 18768 25874 18768 25874 4 _0389_
rlabel metal1 s 3174 24684 3174 24684 4 _0390_
rlabel metal1 s 9200 24922 9200 24922 4 _0391_
rlabel metal1 s 5152 15334 5152 15334 4 _0392_
rlabel metal1 s 7314 26418 7314 26418 4 _0393_
rlabel metal2 s 6854 24888 6854 24888 4 _0394_
rlabel metal1 s 7912 26962 7912 26962 4 _0395_
rlabel metal1 s 2530 10132 2530 10132 4 _0396_
rlabel metal1 s 8878 21658 8878 21658 4 _0397_
rlabel metal2 s 12282 20502 12282 20502 4 _0398_
rlabel metal1 s 11454 21522 11454 21522 4 _0399_
rlabel metal1 s 16238 21522 16238 21522 4 _0400_
rlabel metal1 s 17342 25262 17342 25262 4 _0401_
rlabel metal1 s 13984 19754 13984 19754 4 _0402_
rlabel metal2 s 13018 26214 13018 26214 4 _0403_
rlabel metal1 s 19274 6324 19274 6324 4 _0404_
rlabel metal1 s 3956 22542 3956 22542 4 _0405_
rlabel metal1 s 14536 14382 14536 14382 4 _0406_
rlabel metal1 s 2668 22610 2668 22610 4 _0407_
rlabel metal2 s 2714 21556 2714 21556 4 _0408_
rlabel metal1 s 7314 22202 7314 22202 4 _0409_
rlabel metal1 s 1978 6120 1978 6120 4 _0410_
rlabel metal2 s 8602 20026 8602 20026 4 _0411_
rlabel metal2 s 16882 5372 16882 5372 4 _0412_
rlabel metal1 s 12926 10472 12926 10472 4 _0413_
rlabel metal1 s 20562 6222 20562 6222 4 _0414_
rlabel metal2 s 20194 10795 20194 10795 4 _0415_
rlabel metal1 s 19780 14994 19780 14994 4 _0416_
rlabel metal2 s 6210 13124 6210 13124 4 _0417_
rlabel metal1 s 8188 15130 8188 15130 4 _0418_
rlabel metal2 s 4002 4794 4002 4794 4 _0419_
rlabel metal1 s 1794 6766 1794 6766 4 _0420_
rlabel metal2 s 5934 16252 5934 16252 4 _0421_
rlabel metal2 s 19550 10948 19550 10948 4 _0422_
rlabel metal1 s 12328 11118 12328 11118 4 _0423_
rlabel metal1 s 21436 6426 21436 6426 4 _0424_
rlabel metal1 s 18538 13804 18538 13804 4 _0425_
rlabel metal1 s 19688 12818 19688 12818 4 _0426_
rlabel metal1 s 4738 12614 4738 12614 4 _0427_
rlabel metal2 s 4922 21284 4922 21284 4 _0428_
rlabel metal2 s 4738 4794 4738 4794 4 _0429_
rlabel metal1 s 7360 7514 7360 7514 4 _0430_
rlabel metal1 s 6992 20434 6992 20434 4 _0431_
rlabel metal1 s 15226 20910 15226 20910 4 _0432_
rlabel metal1 s 13478 5202 13478 5202 4 _0433_
rlabel metal1 s 20148 5678 20148 5678 4 _0434_
rlabel metal2 s 6026 23324 6026 23324 4 _0435_
rlabel metal1 s 14214 16524 14214 16524 4 _0436_
rlabel metal1 s 1794 23766 1794 23766 4 _0437_
rlabel metal1 s 5428 23290 5428 23290 4 _0438_
rlabel metal1 s 5612 23834 5612 23834 4 _0439_
rlabel metal2 s 8786 8636 8786 8636 4 _0440_
rlabel metal1 s 6532 19346 6532 19346 4 _0441_
rlabel metal1 s 14628 22610 14628 22610 4 _0442_
rlabel metal1 s 11638 7854 11638 7854 4 _0443_
rlabel metal1 s 5336 25806 5336 25806 4 _0444_
rlabel metal1 s 18124 16082 18124 16082 4 _0445_
rlabel metal1 s 2622 24786 2622 24786 4 _0446_
rlabel metal2 s 4094 25908 4094 25908 4 _0447_
rlabel metal1 s 5060 26010 5060 26010 4 _0448_
rlabel metal1 s 2484 11118 2484 11118 4 _0449_
rlabel metal1 s 9200 18734 9200 18734 4 _0450_
rlabel metal1 s 16652 25738 16652 25738 4 _0451_
rlabel metal1 s 13524 23698 13524 23698 4 _0452_
rlabel metal1 s 21482 7854 21482 7854 4 _0453_
rlabel metal1 s 21666 7922 21666 7922 4 _0454_
rlabel metal2 s 14858 12716 14858 12716 4 _0455_
rlabel metal1 s 14444 12954 14444 12954 4 _0456_
rlabel metal1 s 3680 17850 3680 17850 4 _0457_
rlabel metal2 s 2806 16796 2806 16796 4 _0458_
rlabel metal1 s 8096 10234 8096 10234 4 _0459_
rlabel metal2 s 1886 9724 1886 9724 4 _0460_
rlabel metal1 s 6026 18326 6026 18326 4 _0461_
rlabel metal1 s 15456 11118 15456 11118 4 _0462_
rlabel metal1 s 13202 12410 13202 12410 4 _0463_
rlabel metal1 s 14766 19210 14766 19210 4 _0464_
rlabel metal1 s 18906 12614 18906 12614 4 _0465_
rlabel metal1 s 3818 18734 3818 18734 4 _0466_
rlabel metal2 s 3818 15878 3818 15878 4 _0467_
rlabel metal1 s 7406 5678 7406 5678 4 _0468_
rlabel metal1 s 4048 10030 4048 10030 4 _0469_
rlabel metal1 s 11776 19346 11776 19346 4 _0470_
rlabel metal1 s 18768 9418 18768 9418 4 _0471_
rlabel metal1 s 13892 19482 13892 19482 4 _0472_
rlabel metal1 s 19550 4522 19550 4522 4 _0473_
rlabel metal1 s 14444 19890 14444 19890 4 _0474_
rlabel metal1 s 14536 15674 14536 15674 4 _0475_
rlabel metal1 s 2806 19414 2806 19414 4 _0476_
rlabel metal1 s 2691 20434 2691 20434 4 _0477_
rlabel metal1 s 7774 6970 7774 6970 4 _0478_
rlabel metal1 s 1978 7174 1978 7174 4 _0479_
rlabel metal1 s 11316 16558 11316 16558 4 _0480_
rlabel metal1 s 14214 7276 14214 7276 4 _0481_
rlabel metal1 s 13708 20026 13708 20026 4 _0482_
rlabel metal1 s 7636 23630 7636 23630 4 _0483_
rlabel metal1 s 15548 18258 15548 18258 4 _0484_
rlabel metal1 s 12236 12954 12236 12954 4 _0485_
rlabel metal1 s 6256 24922 6256 24922 4 _0486_
rlabel metal2 s 8786 23290 8786 23290 4 _0487_
rlabel metal1 s 7728 9690 7728 9690 4 _0488_
rlabel metal1 s 7590 18054 7590 18054 4 _0489_
rlabel metal1 s 15548 25262 15548 25262 4 _0490_
rlabel metal2 s 13386 23460 13386 23460 4 _0491_
rlabel metal1 s 17066 13770 17066 13770 4 _0492_
rlabel metal1 s 15916 13294 15916 13294 4 _0493_
rlabel metal1 s 2714 13260 2714 13260 4 _0494_
rlabel metal1 s 3910 14382 3910 14382 4 _0495_
rlabel metal1 s 7452 3026 7452 3026 4 _0496_
rlabel metal1 s 2990 8942 2990 8942 4 _0497_
rlabel metal1 s 5106 3162 5106 3162 4 _0498_
rlabel metal1 s 15548 9554 15548 9554 4 _0499_
rlabel metal1 s 14122 3400 14122 3400 4 _0500_
rlabel metal2 s 16514 7854 16514 7854 4 _0501_
rlabel metal2 s 17526 17340 17526 17340 4 _0502_
rlabel metal1 s 8970 13158 8970 13158 4 _0503_
rlabel metal1 s 5520 17850 5520 17850 4 _0504_
rlabel metal1 s 6716 4114 6716 4114 4 _0505_
rlabel metal1 s 3910 6426 3910 6426 4 _0506_
rlabel metal2 s 11546 16762 11546 16762 4 _0507_
rlabel metal1 s 15870 8058 15870 8058 4 _0508_
rlabel metal2 s 13018 5882 13018 5882 4 _0509_
rlabel metal2 s 21114 4318 21114 4318 4 _0510_
rlabel metal1 s 17710 13770 17710 13770 4 _0511_
rlabel metal2 s 16974 13498 16974 13498 4 _0512_
rlabel metal1 s 3404 12954 3404 12954 4 _0513_
rlabel metal2 s 2806 15470 2806 15470 4 _0514_
rlabel metal1 s 9292 4250 9292 4250 4 _0515_
rlabel metal1 s 4232 8942 4232 8942 4 _0516_
rlabel metal1 s 6256 14994 6256 14994 4 _0517_
rlabel metal2 s 15594 3468 15594 3468 4 _0518_
rlabel metal1 s 13156 4250 13156 4250 4 _0519_
rlabel metal1 s 14674 7888 14674 7888 4 _0520_
rlabel metal1 s 16146 16116 16146 16116 4 _0521_
rlabel metal1 s 9614 11764 9614 11764 4 _0522_
rlabel metal1 s 9292 16082 9292 16082 4 _0523_
rlabel metal2 s 11178 4420 11178 4420 4 _0524_
rlabel metal1 s 9430 7514 9430 7514 4 _0525_
rlabel metal1 s 10396 16218 10396 16218 4 _0526_
rlabel metal1 s 18860 3502 18860 3502 4 _0527_
rlabel metal1 s 13938 7854 13938 7854 4 _0528_
rlabel metal1 s 18308 3910 18308 3910 4 _0529_
rlabel metal1 s 18170 12920 18170 12920 4 _0530_
rlabel metal2 s 6578 12444 6578 12444 4 _0531_
rlabel metal1 s 8648 14586 8648 14586 4 _0532_
rlabel metal2 s 8970 4250 8970 4250 4 _0533_
rlabel metal2 s 6026 9860 6026 9860 4 _0534_
rlabel metal2 s 6394 3638 6394 3638 4 _0535_
rlabel metal2 s 16146 3468 16146 3468 4 _0536_
rlabel metal2 s 13386 3638 13386 3638 4 _0537_
rlabel metal1 s 13754 16082 13754 16082 4 _0538_
rlabel metal2 s 19320 16762 19320 16762 4 _0539_
rlabel metal1 s 10948 13294 10948 13294 4 _0540_
rlabel metal1 s 9476 17850 9476 17850 4 _0541_
rlabel metal2 s 9890 6324 9890 6324 4 _0542_
rlabel metal1 s 10442 9418 10442 9418 4 _0543_
rlabel metal1 s 13202 15980 13202 15980 4 _0544_
rlabel metal2 s 17894 9078 17894 9078 4 _0545_
rlabel metal2 s 13294 7684 13294 7684 4 _0546_
rlabel metal1 s 19412 21386 19412 21386 4 clknet_0_rd_clk
rlabel metal1 s 15088 14790 15088 14790 4 clknet_0_wr_clk
rlabel metal1 s 10902 26010 10902 26010 4 clknet_1_0__leaf_rd_clk
rlabel metal1 s 22310 23154 22310 23154 4 clknet_1_1__leaf_rd_clk
rlabel metal1 s 2162 6766 2162 6766 4 clknet_4_0_0_wr_clk
rlabel metal2 s 21482 3230 21482 3230 4 clknet_4_10_0_wr_clk
rlabel metal2 s 21482 10642 21482 10642 4 clknet_4_11_0_wr_clk
rlabel metal1 s 13478 13362 13478 13362 4 clknet_4_12_0_wr_clk
rlabel metal1 s 14168 21522 14168 21522 4 clknet_4_13_0_wr_clk
rlabel metal1 s 20700 13294 20700 13294 4 clknet_4_14_0_wr_clk
rlabel metal2 s 21574 16354 21574 16354 4 clknet_4_15_0_wr_clk
rlabel metal2 s 2346 12444 2346 12444 4 clknet_4_1_0_wr_clk
rlabel metal2 s 9522 7616 9522 7616 4 clknet_4_2_0_wr_clk
rlabel metal1 s 8786 12274 8786 12274 4 clknet_4_3_0_wr_clk
rlabel metal1 s 2530 18292 2530 18292 4 clknet_4_4_0_wr_clk
rlabel metal1 s 5428 25262 5428 25262 4 clknet_4_5_0_wr_clk
rlabel metal2 s 9706 18530 9706 18530 4 clknet_4_6_0_wr_clk
rlabel metal1 s 8602 23086 8602 23086 4 clknet_4_7_0_wr_clk
rlabel metal1 s 15778 3502 15778 3502 4 clknet_4_8_0_wr_clk
rlabel metal1 s 15778 12614 15778 12614 4 clknet_4_9_0_wr_clk
rlabel metal1 s 20148 26758 20148 26758 4 mem\[0\]\[0\]
rlabel metal1 s 8786 25364 8786 25364 4 mem\[0\]\[1\]
rlabel metal2 s 9338 26112 9338 26112 4 mem\[0\]\[2\]
rlabel metal2 s 8786 26758 8786 26758 4 mem\[0\]\[3\]
rlabel metal1 s 9292 22542 9292 22542 4 mem\[0\]\[4\]
rlabel metal1 s 12558 22202 12558 22202 4 mem\[0\]\[5\]
rlabel metal1 s 17572 26962 17572 26962 4 mem\[0\]\[6\]
rlabel metal2 s 13846 25738 13846 25738 4 mem\[0\]\[7\]
rlabel metal2 s 16514 14212 16514 14212 4 mem\[10\]\[0\]
rlabel metal1 s 4738 13294 4738 13294 4 mem\[10\]\[1\]
rlabel metal1 s 4324 15130 4324 15130 4 mem\[10\]\[2\]
rlabel metal2 s 8234 4386 8234 4386 4 mem\[10\]\[3\]
rlabel metal1 s 3542 10030 3542 10030 4 mem\[10\]\[4\]
rlabel metal1 s 5888 3162 5888 3162 4 mem\[10\]\[5\]
rlabel metal2 s 16238 9792 16238 9792 4 mem\[10\]\[6\]
rlabel metal1 s 13892 3502 13892 3502 4 mem\[10\]\[7\]
rlabel metal1 s 19274 17306 19274 17306 4 mem\[11\]\[0\]
rlabel metal1 s 10074 12614 10074 12614 4 mem\[11\]\[1\]
rlabel metal2 s 5382 19992 5382 19992 4 mem\[11\]\[2\]
rlabel metal1 s 8096 4522 8096 4522 4 mem\[11\]\[3\]
rlabel metal1 s 5336 6630 5336 6630 4 mem\[11\]\[4\]
rlabel metal1 s 13294 17204 13294 17204 4 mem\[11\]\[5\]
rlabel metal2 s 16606 7786 16606 7786 4 mem\[11\]\[6\]
rlabel metal2 s 13386 7191 13386 7191 4 mem\[11\]\[7\]
rlabel metal2 s 18078 13464 18078 13464 4 mem\[12\]\[0\]
rlabel metal1 s 4508 12954 4508 12954 4 mem\[12\]\[1\]
rlabel metal1 s 3542 16082 3542 16082 4 mem\[12\]\[2\]
rlabel metal1 s 10672 3638 10672 3638 4 mem\[12\]\[3\]
rlabel metal1 s 5244 10030 5244 10030 4 mem\[12\]\[4\]
rlabel metal1 s 7176 15674 7176 15674 4 mem\[12\]\[5\]
rlabel metal1 s 16514 4114 16514 4114 4 mem\[12\]\[6\]
rlabel metal1 s 13892 4726 13892 4726 4 mem\[12\]\[7\]
rlabel metal1 s 16928 16490 16928 16490 4 mem\[13\]\[0\]
rlabel metal1 s 10672 12138 10672 12138 4 mem\[13\]\[1\]
rlabel metal2 s 10350 15878 10350 15878 4 mem\[13\]\[2\]
rlabel metal2 s 10258 4182 10258 4182 4 mem\[13\]\[3\]
rlabel metal2 s 10810 7616 10810 7616 4 mem\[13\]\[4\]
rlabel metal1 s 10902 16762 10902 16762 4 mem\[13\]\[5\]
rlabel metal2 s 18354 3264 18354 3264 4 mem\[13\]\[6\]
rlabel metal1 s 14444 8602 14444 8602 4 mem\[13\]\[7\]
rlabel metal1 s 18814 13192 18814 13192 4 mem\[14\]\[0\]
rlabel metal1 s 7544 12886 7544 12886 4 mem\[14\]\[1\]
rlabel metal2 s 9890 15266 9890 15266 4 mem\[14\]\[2\]
rlabel metal2 s 9798 3876 9798 3876 4 mem\[14\]\[3\]
rlabel metal1 s 7222 10710 7222 10710 4 mem\[14\]\[4\]
rlabel metal1 s 6624 3706 6624 3706 4 mem\[14\]\[5\]
rlabel metal1 s 17250 4114 17250 4114 4 mem\[14\]\[6\]
rlabel metal1 s 13892 3706 13892 3706 4 mem\[14\]\[7\]
rlabel metal1 s 19550 16558 19550 16558 4 mem\[15\]\[0\]
rlabel metal1 s 10626 13294 10626 13294 4 mem\[15\]\[1\]
rlabel metal1 s 10074 18394 10074 18394 4 mem\[15\]\[2\]
rlabel metal1 s 10580 6426 10580 6426 4 mem\[15\]\[3\]
rlabel metal1 s 10580 10234 10580 10234 4 mem\[15\]\[4\]
rlabel metal2 s 13570 15878 13570 15878 4 mem\[15\]\[5\]
rlabel metal1 s 17204 9146 17204 9146 4 mem\[15\]\[6\]
rlabel metal1 s 13570 7990 13570 7990 4 mem\[15\]\[7\]
rlabel metal1 s 15226 14314 15226 14314 4 mem\[1\]\[0\]
rlabel metal2 s 3174 22848 3174 22848 4 mem\[1\]\[1\]
rlabel metal1 s 4094 20910 4094 20910 4 mem\[1\]\[2\]
rlabel metal1 s 8418 22576 8418 22576 4 mem\[1\]\[3\]
rlabel metal1 s 4600 6358 4600 6358 4 mem\[1\]\[4\]
rlabel metal2 s 10350 19584 10350 19584 4 mem\[1\]\[5\]
rlabel metal1 s 16468 5338 16468 5338 4 mem\[1\]\[6\]
rlabel metal1 s 13524 10778 13524 10778 4 mem\[1\]\[7\]
rlabel metal1 s 18906 15606 18906 15606 4 mem\[2\]\[0\]
rlabel metal1 s 7038 12954 7038 12954 4 mem\[2\]\[1\]
rlabel metal2 s 7774 14943 7774 14943 4 mem\[2\]\[2\]
rlabel metal2 s 4462 4556 4462 4556 4 mem\[2\]\[3\]
rlabel metal1 s 3496 7446 3496 7446 4 mem\[2\]\[4\]
rlabel metal2 s 7130 16388 7130 16388 4 mem\[2\]\[5\]
rlabel metal1 s 18170 10778 18170 10778 4 mem\[2\]\[6\]
rlabel metal1 s 12926 10234 12926 10234 4 mem\[2\]\[7\]
rlabel metal1 s 19044 14042 19044 14042 4 mem\[3\]\[0\]
rlabel metal1 s 5290 12886 5290 12886 4 mem\[3\]\[1\]
rlabel metal2 s 5658 20944 5658 20944 4 mem\[3\]\[2\]
rlabel metal1 s 5750 4624 5750 4624 4 mem\[3\]\[3\]
rlabel metal1 s 8694 7718 8694 7718 4 mem\[3\]\[4\]
rlabel metal2 s 7406 20672 7406 20672 4 mem\[3\]\[5\]
rlabel metal1 s 15548 21658 15548 21658 4 mem\[3\]\[6\]
rlabel metal1 s 14766 5338 14766 5338 4 mem\[3\]\[7\]
rlabel metal1 s 16008 15946 16008 15946 4 mem\[4\]\[0\]
rlabel metal1 s 4002 23698 4002 23698 4 mem\[4\]\[1\]
rlabel metal2 s 6302 23562 6302 23562 4 mem\[4\]\[2\]
rlabel metal1 s 6256 23562 6256 23562 4 mem\[4\]\[3\]
rlabel metal2 s 10810 8636 10810 8636 4 mem\[4\]\[4\]
rlabel metal1 s 8004 19482 8004 19482 4 mem\[4\]\[5\]
rlabel metal1 s 15364 21998 15364 21998 4 mem\[4\]\[6\]
rlabel metal2 s 12650 7990 12650 7990 4 mem\[4\]\[7\]
rlabel metal2 s 18538 16320 18538 16320 4 mem\[5\]\[0\]
rlabel metal1 s 3404 24038 3404 24038 4 mem\[5\]\[1\]
rlabel metal1 s 5106 25670 5106 25670 4 mem\[5\]\[2\]
rlabel metal1 s 5290 25874 5290 25874 4 mem\[5\]\[3\]
rlabel metal1 s 3818 11730 3818 11730 4 mem\[5\]\[4\]
rlabel metal1 s 10534 18938 10534 18938 4 mem\[5\]\[5\]
rlabel metal1 s 15916 26214 15916 26214 4 mem\[5\]\[6\]
rlabel metal2 s 14306 22984 14306 22984 4 mem\[5\]\[7\]
rlabel metal1 s 15456 13498 15456 13498 4 mem\[6\]\[0\]
rlabel metal1 s 4554 17646 4554 17646 4 mem\[6\]\[1\]
rlabel metal1 s 4094 17238 4094 17238 4 mem\[6\]\[2\]
rlabel metal1 s 8648 10438 8648 10438 4 mem\[6\]\[3\]
rlabel metal2 s 2806 10370 2806 10370 4 mem\[6\]\[4\]
rlabel metal1 s 7958 18734 7958 18734 4 mem\[6\]\[5\]
rlabel metal2 s 16330 10914 16330 10914 4 mem\[6\]\[6\]
rlabel metal1 s 13754 12138 13754 12138 4 mem\[6\]\[7\]
rlabel metal1 s 18952 13430 18952 13430 4 mem\[7\]\[0\]
rlabel metal1 s 4462 18666 4462 18666 4 mem\[7\]\[1\]
rlabel metal1 s 3910 15334 3910 15334 4 mem\[7\]\[2\]
rlabel metal1 s 8372 6426 8372 6426 4 mem\[7\]\[3\]
rlabel metal1 s 5106 9690 5106 9690 4 mem\[7\]\[4\]
rlabel metal1 s 12052 19346 12052 19346 4 mem\[7\]\[5\]
rlabel metal1 s 18078 9894 18078 9894 4 mem\[7\]\[6\]
rlabel metal1 s 14122 19686 14122 19686 4 mem\[7\]\[7\]
rlabel metal1 s 15594 16966 15594 16966 4 mem\[8\]\[0\]
rlabel metal1 s 3358 19890 3358 19890 4 mem\[8\]\[1\]
rlabel metal1 s 3312 20570 3312 20570 4 mem\[8\]\[2\]
rlabel metal1 s 8280 6766 8280 6766 4 mem\[8\]\[3\]
rlabel metal2 s 2806 6698 2806 6698 4 mem\[8\]\[4\]
rlabel metal1 s 13248 16558 13248 16558 4 mem\[8\]\[5\]
rlabel metal2 s 16790 7514 16790 7514 4 mem\[8\]\[6\]
rlabel metal1 s 14260 19822 14260 19822 4 mem\[8\]\[7\]
rlabel metal1 s 16514 18258 16514 18258 4 mem\[9\]\[0\]
rlabel metal1 s 11638 13498 11638 13498 4 mem\[9\]\[1\]
rlabel metal1 s 6670 24854 6670 24854 4 mem\[9\]\[2\]
rlabel metal1 s 7268 23290 7268 23290 4 mem\[9\]\[3\]
rlabel metal1 s 7406 9146 7406 9146 4 mem\[9\]\[4\]
rlabel metal1 s 8188 18258 8188 18258 4 mem\[9\]\[5\]
rlabel metal1 s 16146 25194 16146 25194 4 mem\[9\]\[6\]
rlabel metal2 s 13754 22848 13754 22848 4 mem\[9\]\[7\]
rlabel metal1 s 20838 23018 20838 23018 4 net1
rlabel metal1 s 24932 9690 24932 9690 4 net10
rlabel metal1 s 20792 26418 20792 26418 4 net11
rlabel metal1 s 11776 25126 11776 25126 4 net12
rlabel metal1 s 10350 26928 10350 26928 4 net13
rlabel metal1 s 9706 26010 9706 26010 4 net14
rlabel metal1 s 11408 22542 11408 22542 4 net15
rlabel metal1 s 11822 22712 11822 22712 4 net16
rlabel metal1 s 17618 26418 17618 26418 4 net17
rlabel metal2 s 14490 26588 14490 26588 4 net18
rlabel metal1 s 25806 22610 25806 22610 4 net19
rlabel metal1 s 19550 14484 19550 14484 4 net2
rlabel metal2 s 26358 7327 26358 7327 4 net20
rlabel metal1 s 16560 2346 16560 2346 4 net21
rlabel metal2 s 1518 10234 1518 10234 4 net22
rlabel metal1 s 2162 18258 2162 18258 4 net23
rlabel metal2 s 26450 14586 26450 14586 4 net24
rlabel metal1 s 6256 2346 6256 2346 4 net25
rlabel metal1 s 8878 2414 8878 2414 4 net26
rlabel metal1 s 12972 2414 12972 2414 4 net27
rlabel metal1 s 21436 27438 21436 27438 4 net28
rlabel metal2 s 2070 13124 2070 13124 4 net29
rlabel metal1 s 10488 13158 10488 13158 4 net3
rlabel metal2 s 9798 15164 9798 15164 4 net4
rlabel metal1 s 9246 2516 9246 2516 4 net5
rlabel metal2 s 10166 8466 10166 8466 4 net6
rlabel metal1 s 6164 2618 6164 2618 4 net7
rlabel metal2 s 16422 8738 16422 8738 4 net8
rlabel metal1 s 13478 2482 13478 2482 4 net9
rlabel metal3 s 24449 24956 24449 24956 4 rd_clk
rlabel metal2 s 20102 28509 20102 28509 4 rd_data[0]
rlabel metal1 s 10948 27574 10948 27574 4 rd_data[1]
rlabel metal1 s 10396 27574 10396 27574 4 rd_data[2]
rlabel metal2 s 9798 28509 9798 28509 4 rd_data[3]
rlabel metal2 s 11730 28509 11730 28509 4 rd_data[4]
rlabel metal2 s 12374 28509 12374 28509 4 rd_data[5]
rlabel metal1 s 17480 27574 17480 27574 4 rd_data[6]
rlabel metal2 s 14306 28509 14306 28509 4 rd_data[7]
rlabel metal3 s 26542 22491 26542 22491 4 rd_empty
rlabel metal1 s 20700 27506 20700 27506 4 rd_en
rlabel metal2 s 18906 18496 18906 18496 4 rd_ptr\[0\]
rlabel metal1 s 17434 20536 17434 20536 4 rd_ptr\[1\]
rlabel metal1 s 20010 21488 20010 21488 4 rd_ptr\[2\]
rlabel metal1 s 19274 24786 19274 24786 4 rd_ptr\[3\]
rlabel metal1 s 22816 23698 22816 23698 4 rd_ptr\[4\]
rlabel metal1 s 20424 19686 20424 19686 4 rd_ptr_gray\[0\]
rlabel metal1 s 25162 21488 25162 21488 4 rd_ptr_gray\[1\]
rlabel metal1 s 23322 22678 23322 22678 4 rd_ptr_gray\[2\]
rlabel metal1 s 25208 23494 25208 23494 4 rd_ptr_gray\[3\]
rlabel metal2 s 21758 10268 21758 10268 4 rd_ptr_gray_sync1\[0\]
rlabel metal2 s 25070 14348 25070 14348 4 rd_ptr_gray_sync1\[1\]
rlabel metal2 s 24702 14620 24702 14620 4 rd_ptr_gray_sync1\[2\]
rlabel metal1 s 26128 12886 26128 12886 4 rd_ptr_gray_sync1\[3\]
rlabel metal2 s 22310 14110 22310 14110 4 rd_ptr_gray_sync1\[4\]
rlabel metal1 s 23322 9010 23322 9010 4 rd_ptr_gray_sync2\[0\]
rlabel metal1 s 26174 13158 26174 13158 4 rd_ptr_gray_sync2\[1\]
rlabel metal1 s 25530 14246 25530 14246 4 rd_ptr_gray_sync2\[2\]
rlabel metal1 s 24656 9554 24656 9554 4 rd_ptr_gray_sync2\[3\]
rlabel metal1 s 23644 13838 23644 13838 4 rd_ptr_gray_sync2\[4\]
rlabel metal1 s 22770 25262 22770 25262 4 rd_rst
rlabel metal3 s 1211 26588 1211 26588 4 wr_clk
rlabel metal2 s 25990 14297 25990 14297 4 wr_data[0]
rlabel metal3 s 0 12928 800 13048 4 wr_data[1]
port 17 nsew
rlabel metal3 s 1050 17748 1050 17748 4 wr_data[2]
rlabel metal2 s 8418 1588 8418 1588 4 wr_data[3]
rlabel metal3 s 1050 9588 1050 9588 4 wr_data[4]
rlabel metal2 s 5842 1588 5842 1588 4 wr_data[5]
rlabel metal2 s 16146 1588 16146 1588 4 wr_data[6]
rlabel metal2 s 12926 1027 12926 1027 4 wr_data[7]
rlabel metal1 s 18722 5270 18722 5270 4 wr_en
rlabel metal3 s 26542 7531 26542 7531 4 wr_full
rlabel metal2 s 21390 7174 21390 7174 4 wr_ptr\[0\]
rlabel metal1 s 24288 5678 24288 5678 4 wr_ptr\[1\]
rlabel metal1 s 19228 4590 19228 4590 4 wr_ptr\[2\]
rlabel metal2 s 18538 5746 18538 5746 4 wr_ptr\[3\]
rlabel metal1 s 21022 3434 21022 3434 4 wr_ptr\[4\]
rlabel metal1 s 21344 11866 21344 11866 4 wr_ptr_gray\[0\]
rlabel metal1 s 26128 11322 26128 11322 4 wr_ptr_gray\[1\]
rlabel metal1 s 24748 17578 24748 17578 4 wr_ptr_gray\[2\]
rlabel metal2 s 22310 17663 22310 17663 4 wr_ptr_gray\[3\]
rlabel metal1 s 22586 16422 22586 16422 4 wr_ptr_gray_sync1\[0\]
rlabel metal1 s 24840 17306 24840 17306 4 wr_ptr_gray_sync1\[1\]
rlabel metal2 s 26174 19346 26174 19346 4 wr_ptr_gray_sync1\[2\]
rlabel metal1 s 23460 17850 23460 17850 4 wr_ptr_gray_sync1\[3\]
rlabel metal2 s 22494 17748 22494 17748 4 wr_ptr_gray_sync1\[4\]
rlabel metal2 s 22494 19686 22494 19686 4 wr_ptr_gray_sync2\[0\]
rlabel metal1 s 25944 20366 25944 20366 4 wr_ptr_gray_sync2\[1\]
rlabel metal2 s 24794 21318 24794 21318 4 wr_ptr_gray_sync2\[2\]
rlabel metal1 s 25668 19822 25668 19822 4 wr_ptr_gray_sync2\[3\]
rlabel metal1 s 24058 19822 24058 19822 4 wr_ptr_gray_sync2\[4\]
rlabel metal1 s 26358 10030 26358 10030 4 wr_rst
flabel metal5 s 1056 24716 26912 25116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 20716 26912 21116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 16716 26912 17116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 12716 26912 13116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8716 26912 9116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4716 26912 5116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 23644 2128 24044 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 19644 2128 20044 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 15644 2128 16044 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 11644 2128 12044 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7644 2128 8044 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3644 2128 4044 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 23976 26912 24376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 19976 26912 20376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 15976 26912 16376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 11976 26912 12376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 7976 26912 8376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3976 26912 4376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 22904 2128 23304 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 18904 2128 19304 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 14904 2128 15304 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10904 2128 11304 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 6904 2128 7304 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2904 2128 3304 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 24490 29315 24546 30115 0 FreeSans 280 90 0 0 rd_clk
port 3 nsew
flabel metal2 s 19982 29315 20038 30115 0 FreeSans 280 90 0 0 rd_data[0]
port 4 nsew
flabel metal2 s 10966 29315 11022 30115 0 FreeSans 280 90 0 0 rd_data[1]
port 5 nsew
flabel metal2 s 10322 29315 10378 30115 0 FreeSans 280 90 0 0 rd_data[2]
port 6 nsew
flabel metal2 s 9678 29315 9734 30115 0 FreeSans 280 90 0 0 rd_data[3]
port 7 nsew
flabel metal2 s 11610 29315 11666 30115 0 FreeSans 280 90 0 0 rd_data[4]
port 8 nsew
flabel metal2 s 12254 29315 12310 30115 0 FreeSans 280 90 0 0 rd_data[5]
port 9 nsew
flabel metal2 s 17406 29315 17462 30115 0 FreeSans 280 90 0 0 rd_data[6]
port 10 nsew
flabel metal2 s 14186 29315 14242 30115 0 FreeSans 280 90 0 0 rd_data[7]
port 11 nsew
flabel metal3 s 27171 22448 27971 22568 0 FreeSans 600 0 0 0 rd_empty
port 12 nsew
flabel metal2 s 20626 29315 20682 30115 0 FreeSans 280 90 0 0 rd_en
port 13 nsew
flabel metal2 s 22558 29315 22614 30115 0 FreeSans 280 90 0 0 rd_rst
port 14 nsew
flabel metal3 s 0 26528 800 26648 0 FreeSans 600 0 0 0 wr_clk
port 15 nsew
flabel metal3 s 27171 13608 27971 13728 0 FreeSans 600 0 0 0 wr_data[0]
port 16 nsew
flabel metal3 s 400 12988 400 12988 0 FreeSans 600 0 0 0 wr_data[1]
flabel metal3 s 0 17688 800 17808 0 FreeSans 600 0 0 0 wr_data[2]
port 18 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 wr_data[3]
port 19 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 wr_data[4]
port 20 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 wr_data[5]
port 21 nsew
flabel metal2 s 16118 0 16174 800 0 FreeSans 280 90 0 0 wr_data[6]
port 22 nsew
flabel metal2 s 12898 0 12954 800 0 FreeSans 280 90 0 0 wr_data[7]
port 23 nsew
flabel metal2 s 19338 0 19394 800 0 FreeSans 280 90 0 0 wr_en
port 24 nsew
flabel metal3 s 27171 7488 27971 7608 0 FreeSans 600 0 0 0 wr_full
port 25 nsew
flabel metal3 s 27171 9528 27971 9648 0 FreeSans 600 0 0 0 wr_rst
port 26 nsew
<< properties >>
string FIXED_BBOX 0 0 27971 30115
<< end >>
