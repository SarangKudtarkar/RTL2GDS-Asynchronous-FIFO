magic
tech sky130A
magscale 1 2
timestamp 1756452533
<< nwell >>
rect 1066 2159 26902 27782
<< obsli1 >>
rect 1104 2159 26864 27761
<< obsm1 >>
rect 842 2128 26864 27792
<< metal2 >>
rect 9678 29315 9734 30115
rect 10322 29315 10378 30115
rect 10966 29315 11022 30115
rect 11610 29315 11666 30115
rect 12254 29315 12310 30115
rect 14186 29315 14242 30115
rect 17406 29315 17462 30115
rect 19982 29315 20038 30115
rect 20626 29315 20682 30115
rect 22558 29315 22614 30115
rect 24490 29315 24546 30115
rect 5814 0 5870 800
rect 8390 0 8446 800
rect 12898 0 12954 800
rect 16118 0 16174 800
rect 19338 0 19394 800
<< obsm2 >>
rect 846 29259 9622 29458
rect 9790 29259 10266 29458
rect 10434 29259 10910 29458
rect 11078 29259 11554 29458
rect 11722 29259 12198 29458
rect 12366 29259 14130 29458
rect 14298 29259 17350 29458
rect 17518 29259 19926 29458
rect 20094 29259 20570 29458
rect 20738 29259 22502 29458
rect 22670 29259 24434 29458
rect 24602 29259 26570 29458
rect 846 856 26570 29259
rect 846 800 5758 856
rect 5926 800 8334 856
rect 8502 800 12842 856
rect 13010 800 16062 856
rect 16230 800 19282 856
rect 19450 800 26570 856
<< metal3 >>
rect 0 26528 800 26648
rect 27171 22448 27971 22568
rect 0 17688 800 17808
rect 27171 13608 27971 13728
rect 0 12928 800 13048
rect 0 9528 800 9648
rect 27171 9528 27971 9648
rect 27171 7488 27971 7608
<< obsm3 >>
rect 798 26728 27171 27777
rect 880 26448 27171 26728
rect 798 22648 27171 26448
rect 798 22368 27091 22648
rect 798 17888 27171 22368
rect 880 17608 27171 17888
rect 798 13808 27171 17608
rect 798 13528 27091 13808
rect 798 13128 27171 13528
rect 880 12848 27171 13128
rect 798 9728 27171 12848
rect 880 9448 27091 9728
rect 798 7688 27171 9448
rect 798 7408 27091 7688
rect 798 2143 27171 7408
<< metal4 >>
rect 2904 2128 3304 27792
rect 3644 2128 4044 27792
rect 6904 2128 7304 27792
rect 7644 2128 8044 27792
rect 10904 2128 11304 27792
rect 11644 2128 12044 27792
rect 14904 2128 15304 27792
rect 15644 2128 16044 27792
rect 18904 2128 19304 27792
rect 19644 2128 20044 27792
rect 22904 2128 23304 27792
rect 23644 2128 24044 27792
<< obsm4 >>
rect 5211 6699 6824 26893
rect 7384 6699 7564 26893
rect 8124 6699 10824 26893
rect 11384 6699 11564 26893
rect 12124 6699 14824 26893
rect 15384 6699 15564 26893
rect 16124 6699 18824 26893
rect 19384 6699 19564 26893
rect 20124 6699 22824 26893
rect 23384 6699 23564 26893
rect 24124 6699 24413 26893
<< metal5 >>
rect 1056 24716 26912 25116
rect 1056 23976 26912 24376
rect 1056 20716 26912 21116
rect 1056 19976 26912 20376
rect 1056 16716 26912 17116
rect 1056 15976 26912 16376
rect 1056 12716 26912 13116
rect 1056 11976 26912 12376
rect 1056 8716 26912 9116
rect 1056 7976 26912 8376
rect 1056 4716 26912 5116
rect 1056 3976 26912 4376
<< labels >>
rlabel metal4 s 3644 2128 4044 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7644 2128 8044 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11644 2128 12044 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 15644 2128 16044 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 19644 2128 20044 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 23644 2128 24044 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4716 26912 5116 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8716 26912 9116 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12716 26912 13116 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 16716 26912 17116 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 20716 26912 21116 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 24716 26912 25116 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2904 2128 3304 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6904 2128 7304 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10904 2128 11304 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14904 2128 15304 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 18904 2128 19304 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22904 2128 23304 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3976 26912 4376 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7976 26912 8376 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11976 26912 12376 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 15976 26912 16376 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 19976 26912 20376 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23976 26912 24376 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 24490 29315 24546 30115 6 rd_clk
port 3 nsew signal input
rlabel metal2 s 19982 29315 20038 30115 6 rd_data[0]
port 4 nsew signal output
rlabel metal2 s 10966 29315 11022 30115 6 rd_data[1]
port 5 nsew signal output
rlabel metal2 s 10322 29315 10378 30115 6 rd_data[2]
port 6 nsew signal output
rlabel metal2 s 9678 29315 9734 30115 6 rd_data[3]
port 7 nsew signal output
rlabel metal2 s 11610 29315 11666 30115 6 rd_data[4]
port 8 nsew signal output
rlabel metal2 s 12254 29315 12310 30115 6 rd_data[5]
port 9 nsew signal output
rlabel metal2 s 17406 29315 17462 30115 6 rd_data[6]
port 10 nsew signal output
rlabel metal2 s 14186 29315 14242 30115 6 rd_data[7]
port 11 nsew signal output
rlabel metal3 s 27171 22448 27971 22568 6 rd_empty
port 12 nsew signal output
rlabel metal2 s 20626 29315 20682 30115 6 rd_en
port 13 nsew signal input
rlabel metal2 s 22558 29315 22614 30115 6 rd_rst
port 14 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wr_clk
port 15 nsew signal input
rlabel metal3 s 27171 13608 27971 13728 6 wr_data[0]
port 16 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wr_data[1]
port 17 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wr_data[2]
port 18 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wr_data[3]
port 19 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wr_data[4]
port 20 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wr_data[5]
port 21 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wr_data[6]
port 22 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wr_data[7]
port 23 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wr_en
port 24 nsew signal input
rlabel metal3 s 27171 7488 27971 7608 6 wr_full
port 25 nsew signal output
rlabel metal3 s 27171 9528 27971 9648 6 wr_rst
port 26 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 27971 30115
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2474176
string GDS_FILE /openlane/designs/async_fifo/runs/RUN_2025.08.29_07.26.35/results/signoff/async_fifo.magic.gds
string GDS_START 438888
<< end >>

