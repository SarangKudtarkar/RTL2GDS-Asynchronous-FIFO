VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO async_fifo
  CLASS BLOCK ;
  FOREIGN async_fifo ;
  ORIGIN 0.000 0.000 ;
  SIZE 139.855 BY 150.575 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 18.220 10.640 20.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.220 10.640 40.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.220 10.640 60.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.220 10.640 80.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.220 10.640 100.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.220 10.640 120.220 138.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 23.580 134.560 25.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.580 134.560 45.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 63.580 134.560 65.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 83.580 134.560 85.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 103.580 134.560 105.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 123.580 134.560 125.580 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.520 10.640 16.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.520 10.640 36.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.520 10.640 56.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.520 10.640 76.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.520 10.640 96.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.520 10.640 116.520 138.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.880 134.560 21.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 39.880 134.560 41.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 59.880 134.560 61.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 79.880 134.560 81.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 99.880 134.560 101.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 119.880 134.560 121.880 ;
    END
  END VPWR
  PIN rd_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 146.575 122.730 150.575 ;
    END
  END rd_clk
  PIN rd_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 99.910 146.575 100.190 150.575 ;
    END
  END rd_data[0]
  PIN rd_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 54.830 146.575 55.110 150.575 ;
    END
  END rd_data[1]
  PIN rd_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 51.610 146.575 51.890 150.575 ;
    END
  END rd_data[2]
  PIN rd_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 48.390 146.575 48.670 150.575 ;
    END
  END rd_data[3]
  PIN rd_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 58.050 146.575 58.330 150.575 ;
    END
  END rd_data[4]
  PIN rd_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 61.270 146.575 61.550 150.575 ;
    END
  END rd_data[5]
  PIN rd_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 87.030 146.575 87.310 150.575 ;
    END
  END rd_data[6]
  PIN rd_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 70.930 146.575 71.210 150.575 ;
    END
  END rd_data[7]
  PIN rd_empty
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 135.855 112.240 139.855 112.840 ;
    END
  END rd_empty
  PIN rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 146.575 103.410 150.575 ;
    END
  END rd_en
  PIN rd_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 146.575 113.070 150.575 ;
    END
  END rd_rst
  PIN wr_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wr_clk
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 135.855 68.040 139.855 68.640 ;
    END
  END wr_data[0]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wr_data[1]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wr_data[2]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wr_data[3]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wr_data[4]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wr_data[5]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wr_data[6]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wr_data[7]
  PIN wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wr_en
  PIN wr_full
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 135.855 37.440 139.855 38.040 ;
    END
  END wr_full
  PIN wr_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 135.855 47.640 139.855 48.240 ;
    END
  END wr_rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 134.510 138.910 ;
      LAYER li1 ;
        RECT 5.520 10.795 134.320 138.805 ;
      LAYER met1 ;
        RECT 4.210 10.640 134.320 138.960 ;
      LAYER met2 ;
        RECT 4.230 146.295 48.110 147.290 ;
        RECT 48.950 146.295 51.330 147.290 ;
        RECT 52.170 146.295 54.550 147.290 ;
        RECT 55.390 146.295 57.770 147.290 ;
        RECT 58.610 146.295 60.990 147.290 ;
        RECT 61.830 146.295 70.650 147.290 ;
        RECT 71.490 146.295 86.750 147.290 ;
        RECT 87.590 146.295 99.630 147.290 ;
        RECT 100.470 146.295 102.850 147.290 ;
        RECT 103.690 146.295 112.510 147.290 ;
        RECT 113.350 146.295 122.170 147.290 ;
        RECT 123.010 146.295 132.850 147.290 ;
        RECT 4.230 4.280 132.850 146.295 ;
        RECT 4.230 4.000 28.790 4.280 ;
        RECT 29.630 4.000 41.670 4.280 ;
        RECT 42.510 4.000 64.210 4.280 ;
        RECT 65.050 4.000 80.310 4.280 ;
        RECT 81.150 4.000 96.410 4.280 ;
        RECT 97.250 4.000 132.850 4.280 ;
      LAYER met3 ;
        RECT 3.990 133.640 135.855 138.885 ;
        RECT 4.400 132.240 135.855 133.640 ;
        RECT 3.990 113.240 135.855 132.240 ;
        RECT 3.990 111.840 135.455 113.240 ;
        RECT 3.990 89.440 135.855 111.840 ;
        RECT 4.400 88.040 135.855 89.440 ;
        RECT 3.990 69.040 135.855 88.040 ;
        RECT 3.990 67.640 135.455 69.040 ;
        RECT 3.990 65.640 135.855 67.640 ;
        RECT 4.400 64.240 135.855 65.640 ;
        RECT 3.990 48.640 135.855 64.240 ;
        RECT 4.400 47.240 135.455 48.640 ;
        RECT 3.990 38.440 135.855 47.240 ;
        RECT 3.990 37.040 135.455 38.440 ;
        RECT 3.990 10.715 135.855 37.040 ;
      LAYER met4 ;
        RECT 26.055 33.495 34.120 134.465 ;
        RECT 36.920 33.495 37.820 134.465 ;
        RECT 40.620 33.495 54.120 134.465 ;
        RECT 56.920 33.495 57.820 134.465 ;
        RECT 60.620 33.495 74.120 134.465 ;
        RECT 76.920 33.495 77.820 134.465 ;
        RECT 80.620 33.495 94.120 134.465 ;
        RECT 96.920 33.495 97.820 134.465 ;
        RECT 100.620 33.495 114.120 134.465 ;
        RECT 116.920 33.495 117.820 134.465 ;
        RECT 120.620 33.495 122.065 134.465 ;
  END
END async_fifo
END LIBRARY

