module async_fifo (rd_clk,
    rd_empty,
    rd_en,
    rd_rst,
    wr_clk,
    wr_en,
    wr_full,
    wr_rst,
    rd_data,
    wr_data);
 input rd_clk;
 output rd_empty;
 input rd_en;
 input rd_rst;
 input wr_clk;
 input wr_en;
 output wr_full;
 input wr_rst;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync1[4] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \rd_ptr_gray_sync2[3] ;
 wire \rd_ptr_gray_sync2[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync1[4] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire \wr_ptr_gray_sync2[3] ;
 wire \wr_ptr_gray_sync2[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_wr_clk;
 wire clknet_4_0_0_wr_clk;
 wire clknet_4_1_0_wr_clk;
 wire clknet_4_2_0_wr_clk;
 wire clknet_4_3_0_wr_clk;
 wire clknet_4_4_0_wr_clk;
 wire clknet_4_5_0_wr_clk;
 wire clknet_4_6_0_wr_clk;
 wire clknet_4_7_0_wr_clk;
 wire clknet_4_8_0_wr_clk;
 wire clknet_4_9_0_wr_clk;
 wire clknet_4_10_0_wr_clk;
 wire clknet_4_11_0_wr_clk;
 wire clknet_4_12_0_wr_clk;
 wire clknet_4_13_0_wr_clk;
 wire clknet_4_14_0_wr_clk;
 wire clknet_4_15_0_wr_clk;
 wire clknet_0_rd_clk;
 wire clknet_1_0__leaf_rd_clk;
 wire clknet_1_1__leaf_rd_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;

 sky130_fd_sc_hd__buf_2 _0547_ (.A(\wr_ptr[1] ),
    .X(_0200_));
 sky130_fd_sc_hd__and4_1 _0548_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .C(_0200_),
    .D(\wr_ptr[0] ),
    .X(_0201_));
 sky130_fd_sc_hd__xor2_1 _0549_ (.A(\wr_ptr[4] ),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__a21oi_1 _0550_ (.A1(_0200_),
    .A2(\wr_ptr[0] ),
    .B1(\wr_ptr[2] ),
    .Y(_0203_));
 sky130_fd_sc_hd__xor2_1 _0551_ (.A(\wr_ptr[3] ),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__a2bb2o_1 _0552_ (.A1_N(\rd_ptr_gray_sync2[4] ),
    .A2_N(_0202_),
    .B1(_0204_),
    .B2(\rd_ptr_gray_sync2[2] ),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_4 _0553_ (.A(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__xor2_1 _0554_ (.A(_0200_),
    .B(\wr_ptr[0] ),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _0555_ (.A(\wr_ptr[2] ),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__and3_1 _0556_ (.A(\wr_ptr[2] ),
    .B(_0200_),
    .C(\wr_ptr[0] ),
    .X(_0209_));
 sky130_fd_sc_hd__o21bai_1 _0557_ (.A1(_0203_),
    .A2(_0209_),
    .B1_N(_0207_),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _0558_ (.A(\rd_ptr_gray_sync2[1] ),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_1 _0559_ (.A1(_0208_),
    .A2(_0210_),
    .B1(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _0560_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(_0204_),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _0561_ (.A(\rd_ptr_gray_sync2[3] ),
    .Y(_0214_));
 sky130_fd_sc_hd__a31o_1 _0562_ (.A1(\wr_ptr[2] ),
    .A2(\wr_ptr[1] ),
    .A3(\wr_ptr[0] ),
    .B1(\wr_ptr[3] ),
    .X(_0215_));
 sky130_fd_sc_hd__xnor2_1 _0563_ (.A(\wr_ptr[4] ),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__xnor2_1 _0564_ (.A(_0200_),
    .B(\rd_ptr_gray_sync2[0] ),
    .Y(_0217_));
 sky130_fd_sc_hd__a221o_1 _0565_ (.A1(_0214_),
    .A2(_0216_),
    .B1(_0202_),
    .B2(\rd_ptr_gray_sync2[4] ),
    .C1(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__xor2_1 _0566_ (.A(\wr_ptr[4] ),
    .B(_0215_),
    .X(_0219_));
 sky130_fd_sc_hd__a32o_1 _0567_ (.A1(_0211_),
    .A2(_0208_),
    .A3(_0210_),
    .B1(_0219_),
    .B2(\rd_ptr_gray_sync2[3] ),
    .X(_0220_));
 sky130_fd_sc_hd__or4_1 _0568_ (.A(_0212_),
    .B(_0213_),
    .C(_0218_),
    .D(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_4 _0569_ (.A(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_4 _0570_ (.A(wr_en),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_4 _0571_ (.A(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__o211a_1 _0572_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0224_),
    .C1(_0201_),
    .X(_0225_));
 sky130_fd_sc_hd__xor2_1 _0573_ (.A(\wr_ptr[4] ),
    .B(_0225_),
    .X(_0071_));
 sky130_fd_sc_hd__o21a_2 _0574_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0224_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _0575_ (.A0(\wr_ptr_gray[3] ),
    .A1(_0219_),
    .S(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_1 _0576_ (.A(_0227_),
    .X(_0070_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(_0204_),
    .Y(_0228_));
 sky130_fd_sc_hd__mux2_1 _0578_ (.A0(\wr_ptr_gray[2] ),
    .A1(_0228_),
    .S(_0226_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _0579_ (.A(_0229_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _0580_ (.A(_0208_),
    .B(_0210_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0581_ (.A0(\wr_ptr_gray[1] ),
    .A1(_0230_),
    .S(_0226_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _0582_ (.A(_0231_),
    .X(_0068_));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(_0200_),
    .Y(_0232_));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(\wr_ptr_gray[0] ),
    .A1(_0232_),
    .S(_0226_),
    .X(_0233_));
 sky130_fd_sc_hd__clkbuf_1 _0585_ (.A(_0233_),
    .X(_0067_));
 sky130_fd_sc_hd__o211a_1 _0586_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0224_),
    .C1(_0209_),
    .X(_0234_));
 sky130_fd_sc_hd__o21ba_1 _0587_ (.A1(\wr_ptr[3] ),
    .A2(_0234_),
    .B1_N(_0225_),
    .X(_0066_));
 sky130_fd_sc_hd__nor2_1 _0588_ (.A(_0203_),
    .B(_0209_),
    .Y(_0235_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(\wr_ptr[2] ),
    .A1(_0235_),
    .S(_0226_),
    .X(_0236_));
 sky130_fd_sc_hd__clkbuf_1 _0590_ (.A(_0236_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(_0200_),
    .A1(_0207_),
    .S(_0226_),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_1 _0592_ (.A(_0237_),
    .X(_0064_));
 sky130_fd_sc_hd__xor2_1 _0593_ (.A(\wr_ptr[0] ),
    .B(_0226_),
    .X(_0063_));
 sky130_fd_sc_hd__inv_2 _0594_ (.A(\rd_ptr_gray[1] ),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _0595_ (.A(\wr_ptr_gray_sync2[3] ),
    .Y(_0239_));
 sky130_fd_sc_hd__a22o_1 _0596_ (.A1(_0238_),
    .A2(\wr_ptr_gray_sync2[1] ),
    .B1(_0239_),
    .B2(\rd_ptr_gray[3] ),
    .X(_0240_));
 sky130_fd_sc_hd__xor2_1 _0597_ (.A(\rd_ptr_gray[0] ),
    .B(\wr_ptr_gray_sync2[0] ),
    .X(_0241_));
 sky130_fd_sc_hd__or2b_1 _0598_ (.A(\rd_ptr_gray[3] ),
    .B_N(\wr_ptr_gray_sync2[3] ),
    .X(_0242_));
 sky130_fd_sc_hd__or2b_1 _0599_ (.A(\rd_ptr_gray[2] ),
    .B_N(\wr_ptr_gray_sync2[2] ),
    .X(_0243_));
 sky130_fd_sc_hd__or2b_1 _0600_ (.A(\rd_ptr[4] ),
    .B_N(\wr_ptr_gray_sync2[4] ),
    .X(_0244_));
 sky130_fd_sc_hd__o2111ai_1 _0601_ (.A1(_0238_),
    .A2(\wr_ptr_gray_sync2[1] ),
    .B1(_0242_),
    .C1(_0243_),
    .D1(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _0602_ (.A(\wr_ptr_gray_sync2[2] ),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _0603_ (.A(\wr_ptr_gray_sync2[4] ),
    .Y(_0247_));
 sky130_fd_sc_hd__a22o_1 _0604_ (.A1(\rd_ptr_gray[2] ),
    .A2(_0246_),
    .B1(_0247_),
    .B2(\rd_ptr[4] ),
    .X(_0248_));
 sky130_fd_sc_hd__or4_4 _0605_ (.A(_0240_),
    .B(_0241_),
    .C(_0245_),
    .D(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__and2_1 _0606_ (.A(net1),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__buf_2 _0607_ (.A(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_4 _0608_ (.A(\rd_ptr[3] ),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_4 _0609_ (.A(\rd_ptr[2] ),
    .X(_0253_));
 sky130_fd_sc_hd__and2_1 _0610_ (.A(\rd_ptr[1] ),
    .B(\rd_ptr[0] ),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _0611_ (.A(_0252_),
    .B(_0253_),
    .C(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__clkbuf_4 _0612_ (.A(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_1 _0613_ (.A(_0251_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__xnor2_1 _0614_ (.A(\rd_ptr[4] ),
    .B(_0257_),
    .Y(_0062_));
 sky130_fd_sc_hd__buf_4 _0615_ (.A(\rd_ptr[1] ),
    .X(_0258_));
 sky130_fd_sc_hd__buf_4 _0616_ (.A(\rd_ptr[0] ),
    .X(_0259_));
 sky130_fd_sc_hd__a31o_1 _0617_ (.A1(_0253_),
    .A2(_0258_),
    .A3(_0259_),
    .B1(_0252_),
    .X(_0260_));
 sky130_fd_sc_hd__xor2_1 _0618_ (.A(\rd_ptr[4] ),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(\rd_ptr_gray[3] ),
    .A1(_0261_),
    .S(_0250_),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_1 _0620_ (.A(_0262_),
    .X(_0061_));
 sky130_fd_sc_hd__nor2_1 _0621_ (.A(_0253_),
    .B(_0254_),
    .Y(_0263_));
 sky130_fd_sc_hd__xnor2_1 _0622_ (.A(_0252_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(\rd_ptr_gray[2] ),
    .A1(_0264_),
    .S(_0250_),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _0624_ (.A(_0265_),
    .X(_0060_));
 sky130_fd_sc_hd__or2_2 _0625_ (.A(_0258_),
    .B(_0259_),
    .X(_0266_));
 sky130_fd_sc_hd__xor2_1 _0626_ (.A(_0253_),
    .B(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _0627_ (.A0(\rd_ptr_gray[1] ),
    .A1(_0267_),
    .S(_0250_),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_1 _0628_ (.A(_0268_),
    .X(_0059_));
 sky130_fd_sc_hd__inv_2 _0629_ (.A(_0258_),
    .Y(_0269_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(\rd_ptr_gray[0] ),
    .A1(_0269_),
    .S(_0250_),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _0631_ (.A(_0270_),
    .X(_0058_));
 sky130_fd_sc_hd__and3_1 _0632_ (.A(net1),
    .B(_0249_),
    .C(_0254_),
    .X(_0271_));
 sky130_fd_sc_hd__and2_1 _0633_ (.A(_0253_),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__xor2_1 _0634_ (.A(_0252_),
    .B(_0272_),
    .X(_0057_));
 sky130_fd_sc_hd__nor2_1 _0635_ (.A(_0253_),
    .B(_0271_),
    .Y(_0273_));
 sky130_fd_sc_hd__nor2_1 _0636_ (.A(_0272_),
    .B(_0273_),
    .Y(_0056_));
 sky130_fd_sc_hd__a21oi_1 _0637_ (.A1(_0259_),
    .A2(_0251_),
    .B1(_0258_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor2_1 _0638_ (.A(_0271_),
    .B(_0274_),
    .Y(_0055_));
 sky130_fd_sc_hd__nand2_4 _0639_ (.A(net1),
    .B(_0249_),
    .Y(_0275_));
 sky130_fd_sc_hd__xnor2_1 _0640_ (.A(_0259_),
    .B(_0275_),
    .Y(_0054_));
 sky130_fd_sc_hd__clkbuf_4 _0641_ (.A(\rd_ptr[2] ),
    .X(_0276_));
 sky130_fd_sc_hd__and4b_4 _0642_ (.A_N(_0258_),
    .B(\rd_ptr[0] ),
    .C(_0252_),
    .D(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__and3b_4 _0643_ (.A_N(_0253_),
    .B(_0254_),
    .C(_0252_),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_4 _0644_ (.A(\rd_ptr[3] ),
    .X(_0279_));
 sky130_fd_sc_hd__nor4b_4 _0645_ (.A(_0279_),
    .B(_0258_),
    .C(_0259_),
    .D_N(_0276_),
    .Y(_0280_));
 sky130_fd_sc_hd__a22o_1 _0646_ (.A1(\mem[11][7] ),
    .A2(_0278_),
    .B1(_0280_),
    .B2(\mem[4][7] ),
    .X(_0281_));
 sky130_fd_sc_hd__nor3_4 _0647_ (.A(_0252_),
    .B(_0253_),
    .C(_0266_),
    .Y(_0282_));
 sky130_fd_sc_hd__a211o_1 _0648_ (.A1(\mem[13][7] ),
    .A2(_0277_),
    .B1(_0281_),
    .C1(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__and4bb_4 _0649_ (.A_N(_0279_),
    .B_N(\rd_ptr[0] ),
    .C(\rd_ptr[1] ),
    .D(\rd_ptr[2] ),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _0650_ (.A(\mem[6][7] ),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__nor4b_4 _0651_ (.A(_0279_),
    .B(_0276_),
    .C(_0258_),
    .D_N(\rd_ptr[0] ),
    .Y(_0286_));
 sky130_fd_sc_hd__nor4b_4 _0652_ (.A(_0252_),
    .B(_0253_),
    .C(_0259_),
    .D_N(\rd_ptr[1] ),
    .Y(_0287_));
 sky130_fd_sc_hd__a22o_1 _0653_ (.A1(\mem[1][7] ),
    .A2(_0286_),
    .B1(_0287_),
    .B2(\mem[2][7] ),
    .X(_0288_));
 sky130_fd_sc_hd__and4bb_4 _0654_ (.A_N(_0279_),
    .B_N(_0276_),
    .C(\rd_ptr[1] ),
    .D(\rd_ptr[0] ),
    .X(_0289_));
 sky130_fd_sc_hd__and4bb_4 _0655_ (.A_N(_0258_),
    .B_N(_0259_),
    .C(_0279_),
    .D(\rd_ptr[2] ),
    .X(_0290_));
 sky130_fd_sc_hd__and4b_4 _0656_ (.A_N(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .C(_0276_),
    .D(_0279_),
    .X(_0291_));
 sky130_fd_sc_hd__and4bb_4 _0657_ (.A_N(_0276_),
    .B_N(_0259_),
    .C(\rd_ptr[1] ),
    .D(_0279_),
    .X(_0292_));
 sky130_fd_sc_hd__a22o_1 _0658_ (.A1(\mem[14][7] ),
    .A2(_0291_),
    .B1(_0292_),
    .B2(\mem[10][7] ),
    .X(_0293_));
 sky130_fd_sc_hd__a221o_1 _0659_ (.A1(\mem[3][7] ),
    .A2(_0289_),
    .B1(_0290_),
    .B2(\mem[12][7] ),
    .C1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__and4b_4 _0660_ (.A_N(_0279_),
    .B(_0276_),
    .C(\rd_ptr[1] ),
    .D(\rd_ptr[0] ),
    .X(_0295_));
 sky130_fd_sc_hd__nor4b_4 _0661_ (.A(_0276_),
    .B(_0258_),
    .C(_0259_),
    .D_N(_0279_),
    .Y(_0296_));
 sky130_fd_sc_hd__and4bb_4 _0662_ (.A_N(_0276_),
    .B_N(_0258_),
    .C(\rd_ptr[0] ),
    .D(_0279_),
    .X(_0297_));
 sky130_fd_sc_hd__and4bb_4 _0663_ (.A_N(_0252_),
    .B_N(\rd_ptr[1] ),
    .C(_0259_),
    .D(_0276_),
    .X(_0298_));
 sky130_fd_sc_hd__a22o_1 _0664_ (.A1(\mem[9][7] ),
    .A2(_0297_),
    .B1(_0298_),
    .B2(\mem[5][7] ),
    .X(_0299_));
 sky130_fd_sc_hd__a221o_1 _0665_ (.A1(\mem[7][7] ),
    .A2(_0295_),
    .B1(_0296_),
    .B2(\mem[8][7] ),
    .C1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__or4_1 _0666_ (.A(_0285_),
    .B(_0288_),
    .C(_0294_),
    .D(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__a211o_1 _0667_ (.A1(\mem[15][7] ),
    .A2(_0256_),
    .B1(_0283_),
    .C1(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__or3_4 _0668_ (.A(_0252_),
    .B(_0253_),
    .C(_0266_),
    .X(_0303_));
 sky130_fd_sc_hd__o21a_1 _0669_ (.A1(\mem[0][7] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0304_));
 sky130_fd_sc_hd__a22o_1 _0670_ (.A1(net18),
    .A2(_0275_),
    .B1(_0302_),
    .B2(_0304_),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_1 _0671_ (.A1(\mem[11][6] ),
    .A2(_0278_),
    .B1(_0296_),
    .B2(\mem[8][6] ),
    .X(_0305_));
 sky130_fd_sc_hd__a211o_1 _0672_ (.A1(\mem[15][6] ),
    .A2(_0256_),
    .B1(_0282_),
    .C1(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__a22o_1 _0673_ (.A1(\mem[6][6] ),
    .A2(_0284_),
    .B1(_0292_),
    .B2(\mem[10][6] ),
    .X(_0307_));
 sky130_fd_sc_hd__a22o_1 _0674_ (.A1(\mem[3][6] ),
    .A2(_0289_),
    .B1(_0280_),
    .B2(\mem[4][6] ),
    .X(_0308_));
 sky130_fd_sc_hd__a221o_1 _0675_ (.A1(\mem[9][6] ),
    .A2(_0297_),
    .B1(_0298_),
    .B2(\mem[5][6] ),
    .C1(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__a22o_1 _0676_ (.A1(\mem[13][6] ),
    .A2(_0277_),
    .B1(_0290_),
    .B2(\mem[12][6] ),
    .X(_0310_));
 sky130_fd_sc_hd__a221o_1 _0677_ (.A1(\mem[1][6] ),
    .A2(_0286_),
    .B1(_0291_),
    .B2(\mem[14][6] ),
    .C1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a2111o_1 _0678_ (.A1(\mem[2][6] ),
    .A2(_0287_),
    .B1(_0307_),
    .C1(_0309_),
    .D1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a211o_1 _0679_ (.A1(\mem[7][6] ),
    .A2(_0295_),
    .B1(_0306_),
    .C1(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__o21a_1 _0680_ (.A1(\mem[0][6] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0314_));
 sky130_fd_sc_hd__a22o_1 _0681_ (.A1(net17),
    .A2(_0275_),
    .B1(_0313_),
    .B2(_0314_),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _0682_ (.A1(\mem[15][5] ),
    .A2(_0256_),
    .B1(_0296_),
    .B2(\mem[8][5] ),
    .X(_0315_));
 sky130_fd_sc_hd__a211o_1 _0683_ (.A1(\mem[11][5] ),
    .A2(_0278_),
    .B1(_0315_),
    .C1(_0282_),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _0684_ (.A1(\mem[13][5] ),
    .A2(_0277_),
    .B1(_0298_),
    .B2(\mem[5][5] ),
    .X(_0317_));
 sky130_fd_sc_hd__a22o_1 _0685_ (.A1(\mem[12][5] ),
    .A2(_0290_),
    .B1(_0287_),
    .B2(\mem[2][5] ),
    .X(_0318_));
 sky130_fd_sc_hd__a221o_1 _0686_ (.A1(\mem[9][5] ),
    .A2(_0297_),
    .B1(_0284_),
    .B2(\mem[6][5] ),
    .C1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a22o_1 _0687_ (.A1(\mem[14][5] ),
    .A2(_0291_),
    .B1(_0292_),
    .B2(\mem[10][5] ),
    .X(_0320_));
 sky130_fd_sc_hd__a221o_1 _0688_ (.A1(\mem[3][5] ),
    .A2(_0289_),
    .B1(_0280_),
    .B2(\mem[4][5] ),
    .C1(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__a2111o_1 _0689_ (.A1(\mem[1][5] ),
    .A2(_0286_),
    .B1(_0317_),
    .C1(_0319_),
    .D1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__a211o_1 _0690_ (.A1(\mem[7][5] ),
    .A2(_0295_),
    .B1(_0316_),
    .C1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__o21a_1 _0691_ (.A1(\mem[0][5] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _0692_ (.A1(net16),
    .A2(_0275_),
    .B1(_0323_),
    .B2(_0324_),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_1 _0693_ (.A1(\mem[13][4] ),
    .A2(_0277_),
    .B1(_0289_),
    .B2(\mem[3][4] ),
    .X(_0325_));
 sky130_fd_sc_hd__a211o_1 _0694_ (.A1(\mem[4][4] ),
    .A2(_0280_),
    .B1(_0325_),
    .C1(_0282_),
    .X(_0326_));
 sky130_fd_sc_hd__and2_1 _0695_ (.A(\mem[5][4] ),
    .B(_0298_),
    .X(_0327_));
 sky130_fd_sc_hd__a22o_1 _0696_ (.A1(\mem[14][4] ),
    .A2(_0291_),
    .B1(_0297_),
    .B2(\mem[9][4] ),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _0697_ (.A1(\mem[6][4] ),
    .A2(_0284_),
    .B1(_0292_),
    .B2(\mem[10][4] ),
    .X(_0329_));
 sky130_fd_sc_hd__a221o_1 _0698_ (.A1(\mem[7][4] ),
    .A2(_0295_),
    .B1(_0290_),
    .B2(\mem[12][4] ),
    .C1(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _0699_ (.A1(\mem[8][4] ),
    .A2(_0296_),
    .B1(_0287_),
    .B2(\mem[2][4] ),
    .X(_0331_));
 sky130_fd_sc_hd__a221o_1 _0700_ (.A1(\mem[11][4] ),
    .A2(_0278_),
    .B1(_0286_),
    .B2(\mem[1][4] ),
    .C1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__or4_1 _0701_ (.A(_0327_),
    .B(_0328_),
    .C(_0330_),
    .D(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__a211o_1 _0702_ (.A1(\mem[15][4] ),
    .A2(_0256_),
    .B1(_0326_),
    .C1(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__o21a_1 _0703_ (.A1(\mem[0][4] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _0704_ (.A1(net15),
    .A2(_0275_),
    .B1(_0334_),
    .B2(_0335_),
    .X(_0050_));
 sky130_fd_sc_hd__a22o_1 _0705_ (.A1(\mem[5][3] ),
    .A2(_0298_),
    .B1(_0280_),
    .B2(\mem[4][3] ),
    .X(_0336_));
 sky130_fd_sc_hd__a211o_1 _0706_ (.A1(\mem[6][3] ),
    .A2(_0284_),
    .B1(_0336_),
    .C1(_0282_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _0707_ (.A(\mem[14][3] ),
    .B(_0291_),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _0708_ (.A1(\mem[1][3] ),
    .A2(_0286_),
    .B1(_0297_),
    .B2(\mem[9][3] ),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_1 _0709_ (.A1(\mem[3][3] ),
    .A2(_0289_),
    .B1(_0287_),
    .B2(\mem[2][3] ),
    .X(_0340_));
 sky130_fd_sc_hd__a221o_1 _0710_ (.A1(\mem[11][3] ),
    .A2(_0278_),
    .B1(_0292_),
    .B2(\mem[10][3] ),
    .C1(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _0711_ (.A1(\mem[13][3] ),
    .A2(_0277_),
    .B1(_0290_),
    .B2(\mem[12][3] ),
    .X(_0342_));
 sky130_fd_sc_hd__a221o_1 _0712_ (.A1(\mem[7][3] ),
    .A2(_0295_),
    .B1(_0296_),
    .B2(\mem[8][3] ),
    .C1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__or4_1 _0713_ (.A(_0338_),
    .B(_0339_),
    .C(_0341_),
    .D(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__a211o_1 _0714_ (.A1(\mem[15][3] ),
    .A2(_0256_),
    .B1(_0337_),
    .C1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__o21a_1 _0715_ (.A1(\mem[0][3] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _0716_ (.A1(net14),
    .A2(_0275_),
    .B1(_0345_),
    .B2(_0346_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _0717_ (.A1(\mem[13][2] ),
    .A2(_0277_),
    .B1(_0287_),
    .B2(\mem[2][2] ),
    .X(_0347_));
 sky130_fd_sc_hd__a211o_1 _0718_ (.A1(\mem[14][2] ),
    .A2(_0291_),
    .B1(_0347_),
    .C1(_0282_),
    .X(_0348_));
 sky130_fd_sc_hd__and2_1 _0719_ (.A(\mem[5][2] ),
    .B(_0298_),
    .X(_0349_));
 sky130_fd_sc_hd__a22o_1 _0720_ (.A1(\mem[9][2] ),
    .A2(_0297_),
    .B1(_0280_),
    .B2(\mem[4][2] ),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _0721_ (.A1(\mem[7][2] ),
    .A2(_0295_),
    .B1(_0290_),
    .B2(\mem[12][2] ),
    .X(_0351_));
 sky130_fd_sc_hd__a221o_1 _0722_ (.A1(\mem[6][2] ),
    .A2(_0284_),
    .B1(_0292_),
    .B2(\mem[10][2] ),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _0723_ (.A1(\mem[1][2] ),
    .A2(_0286_),
    .B1(_0296_),
    .B2(\mem[8][2] ),
    .X(_0353_));
 sky130_fd_sc_hd__a221o_1 _0724_ (.A1(\mem[11][2] ),
    .A2(_0278_),
    .B1(_0289_),
    .B2(\mem[3][2] ),
    .C1(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__or4_1 _0725_ (.A(_0349_),
    .B(_0350_),
    .C(_0352_),
    .D(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__a211o_1 _0726_ (.A1(\mem[15][2] ),
    .A2(_0256_),
    .B1(_0348_),
    .C1(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__o21a_1 _0727_ (.A1(\mem[0][2] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_1 _0728_ (.A1(net13),
    .A2(_0275_),
    .B1(_0356_),
    .B2(_0357_),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _0729_ (.A1(\mem[13][1] ),
    .A2(_0277_),
    .B1(_0278_),
    .B2(\mem[11][1] ),
    .X(_0358_));
 sky130_fd_sc_hd__a211o_1 _0730_ (.A1(\mem[9][1] ),
    .A2(_0297_),
    .B1(_0358_),
    .C1(_0282_),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _0731_ (.A(\mem[3][1] ),
    .B(_0289_),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _0732_ (.A1(\mem[14][1] ),
    .A2(_0291_),
    .B1(_0287_),
    .B2(\mem[2][1] ),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _0733_ (.A1(\mem[1][1] ),
    .A2(_0286_),
    .B1(_0298_),
    .B2(\mem[5][1] ),
    .X(_0362_));
 sky130_fd_sc_hd__a221o_1 _0734_ (.A1(\mem[12][1] ),
    .A2(_0290_),
    .B1(_0292_),
    .B2(\mem[10][1] ),
    .C1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__a22o_1 _0735_ (.A1(\mem[4][1] ),
    .A2(_0280_),
    .B1(_0296_),
    .B2(\mem[8][1] ),
    .X(_0364_));
 sky130_fd_sc_hd__a221o_1 _0736_ (.A1(\mem[7][1] ),
    .A2(_0295_),
    .B1(_0284_),
    .B2(\mem[6][1] ),
    .C1(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or4_1 _0737_ (.A(_0360_),
    .B(_0361_),
    .C(_0363_),
    .D(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__a211o_1 _0738_ (.A1(\mem[15][1] ),
    .A2(_0256_),
    .B1(_0359_),
    .C1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__o21a_1 _0739_ (.A1(\mem[0][1] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0368_));
 sky130_fd_sc_hd__a22o_1 _0740_ (.A1(net12),
    .A2(_0275_),
    .B1(_0367_),
    .B2(_0368_),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_1 _0741_ (.A1(\mem[1][0] ),
    .A2(_0286_),
    .B1(_0284_),
    .B2(\mem[6][0] ),
    .X(_0369_));
 sky130_fd_sc_hd__a211o_1 _0742_ (.A1(\mem[10][0] ),
    .A2(_0292_),
    .B1(_0369_),
    .C1(_0282_),
    .X(_0370_));
 sky130_fd_sc_hd__and2_1 _0743_ (.A(\mem[11][0] ),
    .B(_0278_),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_1 _0744_ (.A1(\mem[5][0] ),
    .A2(_0298_),
    .B1(_0287_),
    .B2(\mem[2][0] ),
    .X(_0372_));
 sky130_fd_sc_hd__a22o_1 _0745_ (.A1(\mem[14][0] ),
    .A2(_0291_),
    .B1(_0290_),
    .B2(\mem[12][0] ),
    .X(_0373_));
 sky130_fd_sc_hd__a221o_1 _0746_ (.A1(\mem[7][0] ),
    .A2(_0295_),
    .B1(_0289_),
    .B2(\mem[3][0] ),
    .C1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _0747_ (.A1(\mem[4][0] ),
    .A2(_0280_),
    .B1(_0296_),
    .B2(\mem[8][0] ),
    .X(_0375_));
 sky130_fd_sc_hd__a221o_1 _0748_ (.A1(\mem[13][0] ),
    .A2(_0277_),
    .B1(_0297_),
    .B2(\mem[9][0] ),
    .C1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__or4_1 _0749_ (.A(_0371_),
    .B(_0372_),
    .C(_0374_),
    .D(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__a211o_1 _0750_ (.A1(\mem[15][0] ),
    .A2(_0256_),
    .B1(_0370_),
    .C1(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__o21a_1 _0751_ (.A1(\mem[0][0] ),
    .A2(_0303_),
    .B1(_0251_),
    .X(_0379_));
 sky130_fd_sc_hd__a22o_1 _0752_ (.A1(net11),
    .A2(_0275_),
    .B1(_0378_),
    .B2(_0379_),
    .X(_0046_));
 sky130_fd_sc_hd__nor2_1 _0753_ (.A(_0206_),
    .B(_0222_),
    .Y(net20));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(_0249_),
    .Y(net19));
 sky130_fd_sc_hd__clkbuf_4 _0755_ (.A(rd_rst),
    .X(_0380_));
 sky130_fd_sc_hd__buf_4 _0756_ (.A(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(_0381_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(_0381_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(_0381_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(_0381_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(_0381_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(_0381_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(_0381_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(_0381_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(_0381_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(_0381_),
    .Y(_0009_));
 sky130_fd_sc_hd__buf_4 _0767_ (.A(_0380_),
    .X(_0382_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(_0382_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(_0382_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(_0382_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(_0382_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(_0382_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(_0382_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(_0382_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(_0382_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(_0382_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(_0382_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(_0380_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(_0380_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(net10),
    .Y(_0022_));
 sky130_fd_sc_hd__buf_4 _0781_ (.A(net10),
    .X(_0383_));
 sky130_fd_sc_hd__buf_4 _0782_ (.A(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__inv_2 _0783_ (.A(_0384_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(_0384_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(_0384_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(_0384_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(_0384_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(_0384_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(_0384_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(_0384_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(_0384_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(_0380_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(_0380_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(_0380_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0795_ (.A(_0380_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(_0380_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(_0384_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(_0383_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _0799_ (.A(_0383_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(_0383_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(_0383_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _0802_ (.A(_0383_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(_0383_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(_0383_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(_0383_),
    .Y(_0045_));
 sky130_fd_sc_hd__buf_2 _0806_ (.A(net2),
    .X(_0385_));
 sky130_fd_sc_hd__nor3_2 _0807_ (.A(_0200_),
    .B(\wr_ptr[0] ),
    .C(_0383_),
    .Y(_0386_));
 sky130_fd_sc_hd__nor2_2 _0808_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .Y(_0387_));
 sky130_fd_sc_hd__o2111a_4 _0809_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0386_),
    .C1(_0387_),
    .D1(_0224_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _0810_ (.A0(\mem[0][0] ),
    .A1(_0385_),
    .S(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _0811_ (.A(_0389_),
    .X(_0072_));
 sky130_fd_sc_hd__buf_2 _0812_ (.A(net3),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(\mem[0][1] ),
    .A1(_0390_),
    .S(_0388_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _0814_ (.A(_0391_),
    .X(_0073_));
 sky130_fd_sc_hd__buf_2 _0815_ (.A(net4),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _0816_ (.A0(\mem[0][2] ),
    .A1(_0392_),
    .S(_0388_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0817_ (.A(_0393_),
    .X(_0074_));
 sky130_fd_sc_hd__buf_2 _0818_ (.A(net5),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _0819_ (.A0(\mem[0][3] ),
    .A1(_0394_),
    .S(_0388_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _0820_ (.A(_0395_),
    .X(_0075_));
 sky130_fd_sc_hd__buf_2 _0821_ (.A(net6),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _0822_ (.A0(\mem[0][4] ),
    .A1(_0396_),
    .S(_0388_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _0823_ (.A(_0397_),
    .X(_0076_));
 sky130_fd_sc_hd__buf_2 _0824_ (.A(net7),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(\mem[0][5] ),
    .A1(_0398_),
    .S(_0388_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _0826_ (.A(_0399_),
    .X(_0077_));
 sky130_fd_sc_hd__buf_2 _0827_ (.A(net8),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(\mem[0][6] ),
    .A1(_0400_),
    .S(_0388_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _0829_ (.A(_0401_),
    .X(_0078_));
 sky130_fd_sc_hd__buf_2 _0830_ (.A(net9),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(\mem[0][7] ),
    .A1(_0402_),
    .S(_0388_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _0832_ (.A(_0403_),
    .X(_0079_));
 sky130_fd_sc_hd__and3_2 _0833_ (.A(_0232_),
    .B(\wr_ptr[0] ),
    .C(_0022_),
    .X(_0404_));
 sky130_fd_sc_hd__o2111a_4 _0834_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0387_),
    .C1(_0404_),
    .D1(_0224_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _0835_ (.A0(\mem[1][0] ),
    .A1(_0385_),
    .S(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _0836_ (.A(_0406_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0837_ (.A0(\mem[1][1] ),
    .A1(_0390_),
    .S(_0405_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _0838_ (.A(_0407_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0839_ (.A0(\mem[1][2] ),
    .A1(_0392_),
    .S(_0405_),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_1 _0840_ (.A(_0408_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0841_ (.A0(\mem[1][3] ),
    .A1(_0394_),
    .S(_0405_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _0842_ (.A(_0409_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0843_ (.A0(\mem[1][4] ),
    .A1(_0396_),
    .S(_0405_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _0844_ (.A(_0410_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(\mem[1][5] ),
    .A1(_0398_),
    .S(_0405_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0846_ (.A(_0411_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0847_ (.A0(\mem[1][6] ),
    .A1(_0400_),
    .S(_0405_),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0412_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0849_ (.A0(\mem[1][7] ),
    .A1(_0402_),
    .S(_0405_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _0850_ (.A(_0413_),
    .X(_0087_));
 sky130_fd_sc_hd__and3b_2 _0851_ (.A_N(\wr_ptr[0] ),
    .B(_0022_),
    .C(_0200_),
    .X(_0414_));
 sky130_fd_sc_hd__o2111a_4 _0852_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0387_),
    .C1(_0414_),
    .D1(_0224_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _0853_ (.A0(\mem[2][0] ),
    .A1(_0385_),
    .S(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _0854_ (.A(_0416_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0855_ (.A0(\mem[2][1] ),
    .A1(_0390_),
    .S(_0415_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _0856_ (.A(_0417_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0857_ (.A0(\mem[2][2] ),
    .A1(_0392_),
    .S(_0415_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _0858_ (.A(_0418_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0859_ (.A0(\mem[2][3] ),
    .A1(_0394_),
    .S(_0415_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _0860_ (.A(_0419_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0861_ (.A0(\mem[2][4] ),
    .A1(_0396_),
    .S(_0415_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _0862_ (.A(_0420_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0863_ (.A0(\mem[2][5] ),
    .A1(_0398_),
    .S(_0415_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _0864_ (.A(_0421_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0865_ (.A0(\mem[2][6] ),
    .A1(_0400_),
    .S(_0415_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _0866_ (.A(_0422_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0867_ (.A0(\mem[2][7] ),
    .A1(_0402_),
    .S(_0415_),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _0868_ (.A(_0423_),
    .X(_0095_));
 sky130_fd_sc_hd__and3_1 _0869_ (.A(_0200_),
    .B(\wr_ptr[0] ),
    .C(_0022_),
    .X(_0424_));
 sky130_fd_sc_hd__o2111a_4 _0870_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0387_),
    .C1(_0424_),
    .D1(_0224_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _0871_ (.A0(\mem[3][0] ),
    .A1(_0385_),
    .S(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _0872_ (.A(_0426_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0873_ (.A0(\mem[3][1] ),
    .A1(_0390_),
    .S(_0425_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _0874_ (.A(_0427_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0875_ (.A0(\mem[3][2] ),
    .A1(_0392_),
    .S(_0425_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _0876_ (.A(_0428_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0877_ (.A0(\mem[3][3] ),
    .A1(_0394_),
    .S(_0425_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _0878_ (.A(_0429_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0879_ (.A0(\mem[3][4] ),
    .A1(_0396_),
    .S(_0425_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _0880_ (.A(_0430_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0881_ (.A0(\mem[3][5] ),
    .A1(_0398_),
    .S(_0425_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _0882_ (.A(_0431_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0883_ (.A0(\mem[3][6] ),
    .A1(_0400_),
    .S(_0425_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _0884_ (.A(_0432_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0885_ (.A0(\mem[3][7] ),
    .A1(_0402_),
    .S(_0425_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _0886_ (.A(_0433_),
    .X(_0103_));
 sky130_fd_sc_hd__nor2b_2 _0887_ (.A(\wr_ptr[3] ),
    .B_N(\wr_ptr[2] ),
    .Y(_0434_));
 sky130_fd_sc_hd__o2111a_4 _0888_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0386_),
    .C1(_0434_),
    .D1(_0224_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _0889_ (.A0(\mem[4][0] ),
    .A1(_0385_),
    .S(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _0890_ (.A(_0436_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0891_ (.A0(\mem[4][1] ),
    .A1(_0390_),
    .S(_0435_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _0892_ (.A(_0437_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0893_ (.A0(\mem[4][2] ),
    .A1(_0392_),
    .S(_0435_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _0894_ (.A(_0438_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0895_ (.A0(\mem[4][3] ),
    .A1(_0394_),
    .S(_0435_),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _0896_ (.A(_0439_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0897_ (.A0(\mem[4][4] ),
    .A1(_0396_),
    .S(_0435_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _0898_ (.A(_0440_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0899_ (.A0(\mem[4][5] ),
    .A1(_0398_),
    .S(_0435_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _0900_ (.A(_0441_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0901_ (.A0(\mem[4][6] ),
    .A1(_0400_),
    .S(_0435_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0902_ (.A(_0442_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0903_ (.A0(\mem[4][7] ),
    .A1(_0402_),
    .S(_0435_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _0904_ (.A(_0443_),
    .X(_0111_));
 sky130_fd_sc_hd__o2111a_4 _0905_ (.A1(_0206_),
    .A2(_0222_),
    .B1(_0404_),
    .C1(_0434_),
    .D1(_0224_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(\mem[5][0] ),
    .A1(_0385_),
    .S(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _0907_ (.A(_0445_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0908_ (.A0(\mem[5][1] ),
    .A1(_0390_),
    .S(_0444_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0909_ (.A(_0446_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(\mem[5][2] ),
    .A1(_0392_),
    .S(_0444_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0447_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(\mem[5][3] ),
    .A1(_0394_),
    .S(_0444_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _0913_ (.A(_0448_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(\mem[5][4] ),
    .A1(_0396_),
    .S(_0444_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _0915_ (.A(_0449_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(\mem[5][5] ),
    .A1(_0398_),
    .S(_0444_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _0917_ (.A(_0450_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(\mem[5][6] ),
    .A1(_0400_),
    .S(_0444_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _0919_ (.A(_0451_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(\mem[5][7] ),
    .A1(_0402_),
    .S(_0444_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0452_),
    .X(_0119_));
 sky130_fd_sc_hd__buf_4 _0922_ (.A(_0205_),
    .X(_0453_));
 sky130_fd_sc_hd__buf_4 _0923_ (.A(_0221_),
    .X(_0454_));
 sky130_fd_sc_hd__o2111a_4 _0924_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0414_),
    .C1(_0434_),
    .D1(_0224_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _0925_ (.A0(\mem[6][0] ),
    .A1(_0385_),
    .S(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0926_ (.A(_0456_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0927_ (.A0(\mem[6][1] ),
    .A1(_0390_),
    .S(_0455_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0928_ (.A(_0457_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0929_ (.A0(\mem[6][2] ),
    .A1(_0392_),
    .S(_0455_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0930_ (.A(_0458_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(\mem[6][3] ),
    .A1(_0394_),
    .S(_0455_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _0932_ (.A(_0459_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(\mem[6][4] ),
    .A1(_0396_),
    .S(_0455_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _0934_ (.A(_0460_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(\mem[6][5] ),
    .A1(_0398_),
    .S(_0455_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0936_ (.A(_0461_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(\mem[6][6] ),
    .A1(_0400_),
    .S(_0455_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _0938_ (.A(_0462_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0939_ (.A0(\mem[6][7] ),
    .A1(_0402_),
    .S(_0455_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _0940_ (.A(_0463_),
    .X(_0127_));
 sky130_fd_sc_hd__o2111a_4 _0941_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0424_),
    .C1(_0434_),
    .D1(_0223_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(\mem[7][0] ),
    .A1(_0385_),
    .S(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0943_ (.A(_0465_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(\mem[7][1] ),
    .A1(_0390_),
    .S(_0464_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0945_ (.A(_0466_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(\mem[7][2] ),
    .A1(_0392_),
    .S(_0464_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0947_ (.A(_0467_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(\mem[7][3] ),
    .A1(_0394_),
    .S(_0464_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0468_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(\mem[7][4] ),
    .A1(_0396_),
    .S(_0464_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(_0469_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(\mem[7][5] ),
    .A1(_0398_),
    .S(_0464_),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_1 _0953_ (.A(_0470_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(\mem[7][6] ),
    .A1(_0400_),
    .S(_0464_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0471_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(\mem[7][7] ),
    .A1(_0402_),
    .S(_0464_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _0957_ (.A(_0472_),
    .X(_0135_));
 sky130_fd_sc_hd__nor2b_2 _0958_ (.A(\wr_ptr[2] ),
    .B_N(\wr_ptr[3] ),
    .Y(_0473_));
 sky130_fd_sc_hd__o2111a_4 _0959_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0386_),
    .C1(_0473_),
    .D1(_0223_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(\mem[8][0] ),
    .A1(_0385_),
    .S(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _0961_ (.A(_0475_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(\mem[8][1] ),
    .A1(_0390_),
    .S(_0474_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _0963_ (.A(_0476_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(\mem[8][2] ),
    .A1(_0392_),
    .S(_0474_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_1 _0965_ (.A(_0477_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0966_ (.A0(\mem[8][3] ),
    .A1(_0394_),
    .S(_0474_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _0967_ (.A(_0478_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(\mem[8][4] ),
    .A1(_0396_),
    .S(_0474_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _0969_ (.A(_0479_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(\mem[8][5] ),
    .A1(_0398_),
    .S(_0474_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _0971_ (.A(_0480_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0972_ (.A0(\mem[8][6] ),
    .A1(_0400_),
    .S(_0474_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _0973_ (.A(_0481_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0974_ (.A0(\mem[8][7] ),
    .A1(_0402_),
    .S(_0474_),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _0975_ (.A(_0482_),
    .X(_0143_));
 sky130_fd_sc_hd__o2111a_4 _0976_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0404_),
    .C1(_0473_),
    .D1(_0223_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _0977_ (.A0(\mem[9][0] ),
    .A1(_0385_),
    .S(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _0978_ (.A(_0484_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0979_ (.A0(\mem[9][1] ),
    .A1(_0390_),
    .S(_0483_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(_0485_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0981_ (.A0(\mem[9][2] ),
    .A1(_0392_),
    .S(_0483_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _0982_ (.A(_0486_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0983_ (.A0(\mem[9][3] ),
    .A1(_0394_),
    .S(_0483_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _0984_ (.A(_0487_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0985_ (.A0(\mem[9][4] ),
    .A1(_0396_),
    .S(_0483_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _0986_ (.A(_0488_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0987_ (.A0(\mem[9][5] ),
    .A1(_0398_),
    .S(_0483_),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _0988_ (.A(_0489_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0989_ (.A0(\mem[9][6] ),
    .A1(_0400_),
    .S(_0483_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _0990_ (.A(_0490_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(\mem[9][7] ),
    .A1(_0402_),
    .S(_0483_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(_0491_),
    .X(_0151_));
 sky130_fd_sc_hd__o2111a_4 _0993_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0414_),
    .C1(_0473_),
    .D1(_0223_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(\mem[10][0] ),
    .A1(net2),
    .S(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _0995_ (.A(_0493_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(\mem[10][1] ),
    .A1(net3),
    .S(_0492_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _0997_ (.A(_0494_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(\mem[10][2] ),
    .A1(net4),
    .S(_0492_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(_0495_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(\mem[10][3] ),
    .A1(net5),
    .S(_0492_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(_0496_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(\mem[10][4] ),
    .A1(net6),
    .S(_0492_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(_0497_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(\mem[10][5] ),
    .A1(net7),
    .S(_0492_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _1005_ (.A(_0498_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(\mem[10][6] ),
    .A1(net8),
    .S(_0492_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(_0499_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(\mem[10][7] ),
    .A1(net9),
    .S(_0492_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(_0500_),
    .X(_0159_));
 sky130_fd_sc_hd__o2111a_4 _1010_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0424_),
    .C1(_0473_),
    .D1(_0223_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(\mem[11][0] ),
    .A1(net2),
    .S(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(_0502_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(\mem[11][1] ),
    .A1(net3),
    .S(_0501_),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _1014_ (.A(_0503_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _1015_ (.A0(\mem[11][2] ),
    .A1(net4),
    .S(_0501_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _1016_ (.A(_0504_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _1017_ (.A0(\mem[11][3] ),
    .A1(net5),
    .S(_0501_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _1018_ (.A(_0505_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(\mem[11][4] ),
    .A1(net6),
    .S(_0501_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _1020_ (.A(_0506_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _1021_ (.A0(\mem[11][5] ),
    .A1(net7),
    .S(_0501_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _1022_ (.A(_0507_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(\mem[11][6] ),
    .A1(net8),
    .S(_0501_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _1024_ (.A(_0508_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _1025_ (.A0(\mem[11][7] ),
    .A1(net9),
    .S(_0501_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _1026_ (.A(_0509_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _1027_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .X(_0510_));
 sky130_fd_sc_hd__o2111a_4 _1028_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0386_),
    .C1(_0510_),
    .D1(_0223_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(\mem[12][0] ),
    .A1(net2),
    .S(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(_0512_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(\mem[12][1] ),
    .A1(net3),
    .S(_0511_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_1 _1032_ (.A(_0513_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _1033_ (.A0(\mem[12][2] ),
    .A1(net4),
    .S(_0511_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(_0514_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _1035_ (.A0(\mem[12][3] ),
    .A1(net5),
    .S(_0511_),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(_0515_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _1037_ (.A0(\mem[12][4] ),
    .A1(net6),
    .S(_0511_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(_0516_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(\mem[12][5] ),
    .A1(net7),
    .S(_0511_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _1040_ (.A(_0517_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _1041_ (.A0(\mem[12][6] ),
    .A1(net8),
    .S(_0511_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1042_ (.A(_0518_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _1043_ (.A0(\mem[12][7] ),
    .A1(net9),
    .S(_0511_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_1 _1044_ (.A(_0519_),
    .X(_0175_));
 sky130_fd_sc_hd__o2111a_4 _1045_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0404_),
    .C1(_0510_),
    .D1(_0223_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _1046_ (.A0(\mem[13][0] ),
    .A1(net2),
    .S(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _1047_ (.A(_0521_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _1048_ (.A0(\mem[13][1] ),
    .A1(net3),
    .S(_0520_),
    .X(_0522_));
 sky130_fd_sc_hd__clkbuf_1 _1049_ (.A(_0522_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\mem[13][2] ),
    .A1(net4),
    .S(_0520_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0523_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _1052_ (.A0(\mem[13][3] ),
    .A1(net5),
    .S(_0520_),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_1 _1053_ (.A(_0524_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(\mem[13][4] ),
    .A1(net6),
    .S(_0520_),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _1055_ (.A(_0525_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _1056_ (.A0(\mem[13][5] ),
    .A1(net7),
    .S(_0520_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _1057_ (.A(_0526_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _1058_ (.A0(\mem[13][6] ),
    .A1(net8),
    .S(_0520_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _1059_ (.A(_0527_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _1060_ (.A0(\mem[13][7] ),
    .A1(net9),
    .S(_0520_),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0528_),
    .X(_0183_));
 sky130_fd_sc_hd__o2111a_4 _1062_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0414_),
    .C1(_0510_),
    .D1(_0223_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _1063_ (.A0(\mem[14][0] ),
    .A1(net2),
    .S(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _1064_ (.A(_0530_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _1065_ (.A0(\mem[14][1] ),
    .A1(net3),
    .S(_0529_),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _1066_ (.A(_0531_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _1067_ (.A0(\mem[14][2] ),
    .A1(net4),
    .S(_0529_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1068_ (.A(_0532_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _1069_ (.A0(\mem[14][3] ),
    .A1(net5),
    .S(_0529_),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_1 _1070_ (.A(_0533_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _1071_ (.A0(\mem[14][4] ),
    .A1(net6),
    .S(_0529_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_1 _1072_ (.A(_0534_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _1073_ (.A0(\mem[14][5] ),
    .A1(net7),
    .S(_0529_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _1074_ (.A(_0535_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _1075_ (.A0(\mem[14][6] ),
    .A1(net8),
    .S(_0529_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1076_ (.A(_0536_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _1077_ (.A0(\mem[14][7] ),
    .A1(net9),
    .S(_0529_),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _1078_ (.A(_0537_),
    .X(_0191_));
 sky130_fd_sc_hd__o2111a_4 _1079_ (.A1(_0453_),
    .A2(_0454_),
    .B1(_0223_),
    .C1(_0022_),
    .D1(_0201_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _1080_ (.A0(\mem[15][0] ),
    .A1(net2),
    .S(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _1081_ (.A(_0539_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _1082_ (.A0(\mem[15][1] ),
    .A1(net3),
    .S(_0538_),
    .X(_0540_));
 sky130_fd_sc_hd__clkbuf_1 _1083_ (.A(_0540_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _1084_ (.A0(\mem[15][2] ),
    .A1(net4),
    .S(_0538_),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_1 _1085_ (.A(_0541_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _1086_ (.A0(\mem[15][3] ),
    .A1(net5),
    .S(_0538_),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_1 _1087_ (.A(_0542_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _1088_ (.A0(\mem[15][4] ),
    .A1(net6),
    .S(_0538_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _1089_ (.A(_0543_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(\mem[15][5] ),
    .A1(net7),
    .S(_0538_),
    .X(_0544_));
 sky130_fd_sc_hd__clkbuf_1 _1091_ (.A(_0544_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _1092_ (.A0(\mem[15][6] ),
    .A1(net8),
    .S(_0538_),
    .X(_0545_));
 sky130_fd_sc_hd__clkbuf_1 _1093_ (.A(_0545_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _1094_ (.A0(\mem[15][7] ),
    .A1(net9),
    .S(_0538_),
    .X(_0546_));
 sky130_fd_sc_hd__clkbuf_1 _1095_ (.A(_0546_),
    .X(_0199_));
 sky130_fd_sc_hd__dfrtp_1 _1096_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray[0] ),
    .RESET_B(_0000_),
    .Q(\wr_ptr_gray_sync1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray[1] ),
    .RESET_B(_0001_),
    .Q(\wr_ptr_gray_sync1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray[2] ),
    .RESET_B(_0002_),
    .Q(\wr_ptr_gray_sync1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1099_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray[3] ),
    .RESET_B(_0003_),
    .Q(\wr_ptr_gray_sync1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1100_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr[4] ),
    .RESET_B(_0004_),
    .Q(\wr_ptr_gray_sync1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1101_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray_sync1[0] ),
    .RESET_B(_0005_),
    .Q(\wr_ptr_gray_sync2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray_sync1[1] ),
    .RESET_B(_0006_),
    .Q(\wr_ptr_gray_sync2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray_sync1[2] ),
    .RESET_B(_0007_),
    .Q(\wr_ptr_gray_sync2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray_sync1[3] ),
    .RESET_B(_0008_),
    .Q(\wr_ptr_gray_sync2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(\wr_ptr_gray_sync1[4] ),
    .RESET_B(_0009_),
    .Q(\wr_ptr_gray_sync2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0046_),
    .RESET_B(_0010_),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_1 _1107_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0047_),
    .RESET_B(_0011_),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0048_),
    .RESET_B(_0012_),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0049_),
    .RESET_B(_0013_),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0050_),
    .RESET_B(_0014_),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0051_),
    .RESET_B(_0015_),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0052_),
    .RESET_B(_0016_),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0053_),
    .RESET_B(_0017_),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_4 _1114_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0054_),
    .RESET_B(_0018_),
    .Q(\rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1115_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0055_),
    .RESET_B(_0019_),
    .Q(\rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1116_ (.CLK(clknet_1_0__leaf_rd_clk),
    .D(_0056_),
    .RESET_B(_0020_),
    .Q(\rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1117_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(_0057_),
    .RESET_B(_0021_),
    .Q(\rd_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(clknet_4_11_0_wr_clk),
    .D(\rd_ptr_gray[0] ),
    .RESET_B(_0022_),
    .Q(\rd_ptr_gray_sync1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_4_15_0_wr_clk),
    .D(\rd_ptr_gray[1] ),
    .RESET_B(_0023_),
    .Q(\rd_ptr_gray_sync1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_4_14_0_wr_clk),
    .D(\rd_ptr_gray[2] ),
    .RESET_B(_0024_),
    .Q(\rd_ptr_gray_sync1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1121_ (.CLK(clknet_4_15_0_wr_clk),
    .D(\rd_ptr_gray[3] ),
    .RESET_B(_0025_),
    .Q(\rd_ptr_gray_sync1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1122_ (.CLK(clknet_4_15_0_wr_clk),
    .D(\rd_ptr[4] ),
    .RESET_B(_0026_),
    .Q(\rd_ptr_gray_sync1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1123_ (.CLK(clknet_4_11_0_wr_clk),
    .D(\rd_ptr_gray_sync1[0] ),
    .RESET_B(_0027_),
    .Q(\rd_ptr_gray_sync2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1124_ (.CLK(clknet_4_14_0_wr_clk),
    .D(\rd_ptr_gray_sync1[1] ),
    .RESET_B(_0028_),
    .Q(\rd_ptr_gray_sync2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_4_15_0_wr_clk),
    .D(\rd_ptr_gray_sync1[2] ),
    .RESET_B(_0029_),
    .Q(\rd_ptr_gray_sync2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_4_15_0_wr_clk),
    .D(\rd_ptr_gray_sync1[3] ),
    .RESET_B(_0030_),
    .Q(\rd_ptr_gray_sync2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_4_14_0_wr_clk),
    .D(\rd_ptr_gray_sync1[4] ),
    .RESET_B(_0031_),
    .Q(\rd_ptr_gray_sync2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(_0058_),
    .RESET_B(_0032_),
    .Q(\rd_ptr_gray[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(_0059_),
    .RESET_B(_0033_),
    .Q(\rd_ptr_gray[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(_0060_),
    .RESET_B(_0034_),
    .Q(\rd_ptr_gray[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(_0061_),
    .RESET_B(_0035_),
    .Q(\rd_ptr_gray[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1132_ (.CLK(clknet_1_1__leaf_rd_clk),
    .D(_0062_),
    .RESET_B(_0036_),
    .Q(\rd_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1133_ (.CLK(clknet_4_10_0_wr_clk),
    .D(_0063_),
    .RESET_B(_0037_),
    .Q(\wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_4_10_0_wr_clk),
    .D(_0064_),
    .RESET_B(_0038_),
    .Q(\wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1135_ (.CLK(clknet_4_10_0_wr_clk),
    .D(_0065_),
    .RESET_B(_0039_),
    .Q(\wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1136_ (.CLK(clknet_4_10_0_wr_clk),
    .D(_0066_),
    .RESET_B(_0040_),
    .Q(\wr_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(clknet_4_11_0_wr_clk),
    .D(_0067_),
    .RESET_B(_0041_),
    .Q(\wr_ptr_gray[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(clknet_4_11_0_wr_clk),
    .D(_0068_),
    .RESET_B(_0042_),
    .Q(\wr_ptr_gray[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(clknet_4_11_0_wr_clk),
    .D(_0069_),
    .RESET_B(_0043_),
    .Q(\wr_ptr_gray[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1140_ (.CLK(clknet_4_14_0_wr_clk),
    .D(_0070_),
    .RESET_B(_0044_),
    .Q(\wr_ptr_gray[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1141_ (.CLK(clknet_4_10_0_wr_clk),
    .D(_0071_),
    .RESET_B(_0045_),
    .Q(\wr_ptr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(clknet_4_13_0_wr_clk),
    .D(_0072_),
    .Q(\mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0073_),
    .Q(\mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0074_),
    .Q(\mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1145_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0075_),
    .Q(\mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0076_),
    .Q(\mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0077_),
    .Q(\mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.CLK(clknet_4_13_0_wr_clk),
    .D(_0078_),
    .Q(\mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0079_),
    .Q(\mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0080_),
    .Q(\mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0081_),
    .Q(\mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0082_),
    .Q(\mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0083_),
    .Q(\mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0084_),
    .Q(\mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0085_),
    .Q(\mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.CLK(clknet_4_8_0_wr_clk),
    .D(_0086_),
    .Q(\mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.CLK(clknet_4_9_0_wr_clk),
    .D(_0087_),
    .Q(\mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1158_ (.CLK(clknet_4_15_0_wr_clk),
    .D(_0088_),
    .Q(\mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0089_),
    .Q(\mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0090_),
    .Q(\mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0091_),
    .Q(\mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0092_),
    .Q(\mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0093_),
    .Q(\mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.CLK(clknet_4_11_0_wr_clk),
    .D(_0094_),
    .Q(\mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.CLK(clknet_4_3_0_wr_clk),
    .D(_0095_),
    .Q(\mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.CLK(clknet_4_14_0_wr_clk),
    .D(_0096_),
    .Q(\mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0097_),
    .Q(\mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0098_),
    .Q(\mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0099_),
    .Q(\mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1170_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0100_),
    .Q(\mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0101_),
    .Q(\mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1172_ (.CLK(clknet_4_13_0_wr_clk),
    .D(_0102_),
    .Q(\mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1173_ (.CLK(clknet_4_8_0_wr_clk),
    .D(_0103_),
    .Q(\mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1174_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0104_),
    .Q(\mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0105_),
    .Q(\mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1176_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0106_),
    .Q(\mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1177_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0107_),
    .Q(\mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1178_ (.CLK(clknet_4_3_0_wr_clk),
    .D(_0108_),
    .Q(\mem[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0109_),
    .Q(\mem[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.CLK(clknet_4_13_0_wr_clk),
    .D(_0110_),
    .Q(\mem[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0111_),
    .Q(\mem[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0112_),
    .Q(\mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0113_),
    .Q(\mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0114_),
    .Q(\mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0115_),
    .Q(\mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1186_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0116_),
    .Q(\mem[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0117_),
    .Q(\mem[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1188_ (.CLK(clknet_4_13_0_wr_clk),
    .D(_0118_),
    .Q(\mem[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0119_),
    .Q(\mem[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1190_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0120_),
    .Q(\mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1191_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0121_),
    .Q(\mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0122_),
    .Q(\mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.CLK(clknet_4_3_0_wr_clk),
    .D(_0123_),
    .Q(\mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1194_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0124_),
    .Q(\mem[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0125_),
    .Q(\mem[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1196_ (.CLK(clknet_4_9_0_wr_clk),
    .D(_0126_),
    .Q(\mem[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.CLK(clknet_4_9_0_wr_clk),
    .D(_0127_),
    .Q(\mem[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1198_ (.CLK(clknet_4_14_0_wr_clk),
    .D(_0128_),
    .Q(\mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1199_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0129_),
    .Q(\mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1200_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0130_),
    .Q(\mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0131_),
    .Q(\mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0132_),
    .Q(\mem[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1203_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0133_),
    .Q(\mem[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1204_ (.CLK(clknet_4_11_0_wr_clk),
    .D(_0134_),
    .Q(\mem[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0135_),
    .Q(\mem[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1206_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0136_),
    .Q(\mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1207_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0137_),
    .Q(\mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0138_),
    .Q(\mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1209_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0139_),
    .Q(\mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1210_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0140_),
    .Q(\mem[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1211_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0141_),
    .Q(\mem[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1212_ (.CLK(clknet_4_8_0_wr_clk),
    .D(_0142_),
    .Q(\mem[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0143_),
    .Q(\mem[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1214_ (.CLK(clknet_4_13_0_wr_clk),
    .D(_0144_),
    .Q(\mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0145_),
    .Q(\mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.CLK(clknet_4_5_0_wr_clk),
    .D(_0146_),
    .Q(\mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0147_),
    .Q(\mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0148_),
    .Q(\mem[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1219_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0149_),
    .Q(\mem[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1220_ (.CLK(clknet_4_13_0_wr_clk),
    .D(_0150_),
    .Q(\mem[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1221_ (.CLK(clknet_4_7_0_wr_clk),
    .D(_0151_),
    .Q(\mem[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1222_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0152_),
    .Q(\mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1223_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0153_),
    .Q(\mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1224_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0154_),
    .Q(\mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1225_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0155_),
    .Q(\mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1226_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0156_),
    .Q(\mem[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1227_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0157_),
    .Q(\mem[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1228_ (.CLK(clknet_4_9_0_wr_clk),
    .D(_0158_),
    .Q(\mem[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1229_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0159_),
    .Q(\mem[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1230_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0160_),
    .Q(\mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1231_ (.CLK(clknet_4_3_0_wr_clk),
    .D(_0161_),
    .Q(\mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1232_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0162_),
    .Q(\mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1233_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0163_),
    .Q(\mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0164_),
    .Q(\mem[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0165_),
    .Q(\mem[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1236_ (.CLK(clknet_4_8_0_wr_clk),
    .D(_0166_),
    .Q(\mem[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0167_),
    .Q(\mem[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1238_ (.CLK(clknet_4_9_0_wr_clk),
    .D(_0168_),
    .Q(\mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1239_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0169_),
    .Q(\mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0170_),
    .Q(\mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0171_),
    .Q(\mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0172_),
    .Q(\mem[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_4_4_0_wr_clk),
    .D(_0173_),
    .Q(\mem[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1244_ (.CLK(clknet_4_8_0_wr_clk),
    .D(_0174_),
    .Q(\mem[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1245_ (.CLK(clknet_4_8_0_wr_clk),
    .D(_0175_),
    .Q(\mem[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0176_),
    .Q(\mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_4_3_0_wr_clk),
    .D(_0177_),
    .Q(\mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0178_),
    .Q(\mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0179_),
    .Q(\mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_4_3_0_wr_clk),
    .D(_0180_),
    .Q(\mem[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0181_),
    .Q(\mem[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_4_10_0_wr_clk),
    .D(_0182_),
    .Q(\mem[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_4_9_0_wr_clk),
    .D(_0183_),
    .Q(\mem[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_4_12_0_wr_clk),
    .D(_0184_),
    .Q(\mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0185_),
    .Q(\mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0186_),
    .Q(\mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1257_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0187_),
    .Q(\mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_4_1_0_wr_clk),
    .D(_0188_),
    .Q(\mem[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1259_ (.CLK(clknet_4_0_0_wr_clk),
    .D(_0189_),
    .Q(\mem[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_4_8_0_wr_clk),
    .D(_0190_),
    .Q(\mem[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0191_),
    .Q(\mem[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_4_15_0_wr_clk),
    .D(_0192_),
    .Q(\mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_4_9_0_wr_clk),
    .D(_0193_),
    .Q(\mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0194_),
    .Q(\mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0195_),
    .Q(\mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_4_3_0_wr_clk),
    .D(_0196_),
    .Q(\mem[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_4_6_0_wr_clk),
    .D(_0197_),
    .Q(\mem[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_4_11_0_wr_clk),
    .D(_0198_),
    .Q(\mem[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_4_2_0_wr_clk),
    .D(_0199_),
    .Q(\mem[15][7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_313 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(net28),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(net24),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(net29),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(net23),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(net26),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(net22),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(net25),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(net21),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(net27),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(wr_rst),
    .X(net10));
 sky130_fd_sc_hd__buf_1 output11 (.A(net11),
    .X(rd_data[0]));
 sky130_fd_sc_hd__buf_1 output12 (.A(net12),
    .X(rd_data[1]));
 sky130_fd_sc_hd__buf_1 output13 (.A(net13),
    .X(rd_data[2]));
 sky130_fd_sc_hd__buf_1 output14 (.A(net14),
    .X(rd_data[3]));
 sky130_fd_sc_hd__buf_1 output15 (.A(net15),
    .X(rd_data[4]));
 sky130_fd_sc_hd__buf_1 output16 (.A(net16),
    .X(rd_data[5]));
 sky130_fd_sc_hd__buf_1 output17 (.A(net17),
    .X(rd_data[6]));
 sky130_fd_sc_hd__buf_1 output18 (.A(net18),
    .X(rd_data[7]));
 sky130_fd_sc_hd__buf_1 output19 (.A(net19),
    .X(rd_empty));
 sky130_fd_sc_hd__buf_1 output20 (.A(net20),
    .X(wr_full));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wr_clk (.A(wr_clk),
    .X(clknet_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_0_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_1_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_2_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_3_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_4_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_5_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_6_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_7_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_8_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_9_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_10_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_11_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_12_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_13_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_14_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wr_clk (.A(clknet_0_wr_clk),
    .X(clknet_4_15_0_wr_clk));
 sky130_fd_sc_hd__clkinv_1 clkload0 (.A(clknet_4_0_0_wr_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_4_1_0_wr_clk));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_4_2_0_wr_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_4_3_0_wr_clk));
 sky130_fd_sc_hd__bufinv_16 clkload4 (.A(clknet_4_4_0_wr_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_4_6_0_wr_clk));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_4_7_0_wr_clk));
 sky130_fd_sc_hd__inv_6 clkload7 (.A(clknet_4_8_0_wr_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_4_9_0_wr_clk));
 sky130_fd_sc_hd__inv_8 clkload9 (.A(clknet_4_10_0_wr_clk));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_4_11_0_wr_clk));
 sky130_fd_sc_hd__clkinv_4 clkload11 (.A(clknet_4_12_0_wr_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_4_13_0_wr_clk));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_4_14_0_wr_clk));
 sky130_fd_sc_hd__inv_6 clkload14 (.A(clknet_4_15_0_wr_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_rd_clk (.A(rd_clk),
    .X(clknet_0_rd_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_rd_clk (.A(clknet_0_rd_clk),
    .X(clknet_1_0__leaf_rd_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_rd_clk (.A(clknet_0_rd_clk),
    .X(clknet_1_1__leaf_rd_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload15 (.A(clknet_1_0__leaf_rd_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(wr_data[6]),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(wr_data[4]),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(wr_data[2]),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(wr_data[0]),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(wr_data[5]),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(wr_data[3]),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(wr_data[7]),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(rd_en),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(wr_data[1]),
    .X(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(wr_data[0]));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
endmodule
